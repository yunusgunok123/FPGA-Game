
module main(
input wire CLK,             	// 25.175 MHz clock
input wire RESET,             	// Reset signal
input wire Weapon_switch, 		// To switch the current weapon (Button3)
input wire Fire, 		// Fire button (Button4)
input wire Rotate_CW, 			// To rotate 22.5 degrees in clockwise direction (Button2)
input wire Rotate_CCW, 			// To rotate 22.5 degrees in counter-clockwise direction (Button1)
input wire Interaction,		    // Used as an interaction button for "Try again", "OKAY" (Button5)
output wire hsync,              // Horizontal sync output
output wire vsync,              // Vertical sync output
output wire[7:0] red,		    // Pixel color information about red color
output wire[7:0] green,		    // Pixel color information about green color
output wire[7:0] blue,		    // Pixel color information about blue color
output reg Alive					// Player is alive or not
);

wire[9:0] hc;
wire[9:0] vc;
wire is_blanking;

VGA_init(.CLK(CLK),.RESET(RESET),.hsync(hsync),.vsync(vsync),.hc(hc),.vc(vc),.is_blanking(is_blanking));

parameter [23:0] color0  = {8'd026, 8'd028, 8'd043};
parameter [23:0] color1  = {8'd093, 8'd038, 8'd093};
parameter [23:0] color2  = {8'd178, 8'd062, 8'd083};
parameter [23:0] color3  = {8'd239, 8'd125, 8'd088};
parameter [23:0] color4  = {8'd255, 8'd205, 8'd118};
parameter [23:0] color5  = {8'd168, 8'd240, 8'd112};
parameter [23:0] color6  = {8'd054, 8'd184, 8'd101};
parameter [23:0] color7  = {8'd036, 8'd113, 8'd121};
parameter [23:0] color8  = {8'd042, 8'd054, 8'd112};
parameter [23:0] color9  = {8'd059, 8'd093, 8'd201};
parameter [23:0] color10 = {8'd065, 8'd166, 8'd246};
parameter [23:0] color11 = {8'd115, 8'd239, 8'd247};
parameter [23:0] color12 = {8'd244, 8'd244, 8'd244};
parameter [23:0] color13 = {8'd149, 8'd176, 8'd195};
parameter [23:0] color14 = {8'd086, 8'd107, 8'd134};
parameter [23:0] color15 = {8'd050, 8'd060, 8'd087};

reg[3:0] pixel;

assign red = (is_blanking) ? 8'b00000000:
	(pixel == 4'd0) ? color0[23:16]:
	(pixel == 4'd1) ? color1[23:16]:
	(pixel == 4'd2) ? color2[23:16]:
	(pixel == 4'd3) ? color3[23:16]:
	(pixel == 4'd4) ? color4[23:16]:
	(pixel == 4'd5) ? color5[23:16]:
	(pixel == 4'd6) ? color6[23:16]:
	(pixel == 4'd7) ? color7[23:16]:
	(pixel == 4'd8) ? color8[23:16]:
	(pixel == 4'd9) ? color9[23:16]:
	(pixel == 4'd10) ? color10[23:16]:
	(pixel == 4'd11) ? color11[23:16]:
	(pixel == 4'd12) ? color12[23:16]:
	(pixel == 4'd13) ? color13[23:16]:
	(pixel == 4'd14) ? color14[23:16]:
	color15[23:16];

assign green = (is_blanking) ? 8'b00000000:
	(pixel == 4'd0) ? color0[15:8]:
	(pixel == 4'd1) ? color1[15:8]:
	(pixel == 4'd2) ? color2[15:8]:
	(pixel == 4'd3) ? color3[15:8]:
	(pixel == 4'd4) ? color4[15:8]:
	(pixel == 4'd5) ? color5[15:8]:
	(pixel == 4'd6) ? color6[15:8]:
	(pixel == 4'd7) ? color7[15:8]:
	(pixel == 4'd8) ? color8[15:8]:
	(pixel == 4'd9) ? color9[15:8]:
	(pixel == 4'd10) ? color10[15:8]:
	(pixel == 4'd11) ? color11[15:8]:
	(pixel == 4'd12) ? color12[15:8]:
	(pixel == 4'd13) ? color13[15:8]:
	(pixel == 4'd14) ? color14[15:8]:
	color15[15:8];

assign blue = (is_blanking) ? 8'b00000000:
	(pixel == 4'd0) ? color0[7:0]:
	(pixel == 4'd1) ? color1[7:0]:
	(pixel == 4'd2) ? color2[7:0]:
	(pixel == 4'd3) ? color3[7:0]:
	(pixel == 4'd4) ? color4[7:0]:
	(pixel == 4'd5) ? color5[7:0]:
	(pixel == 4'd6) ? color6[7:0]:
	(pixel == 4'd7) ? color7[7:0]:
	(pixel == 4'd8) ? color8[7:0]:
	(pixel == 4'd9) ? color9[7:0]:
	(pixel == 4'd10) ? color10[7:0]:
	(pixel == 4'd11) ? color11[7:0]:
	(pixel == 4'd12) ? color12[7:0]:
	(pixel == 4'd13) ? color13[7:0]:
	(pixel == 4'd14) ? color14[7:0]:
	color15[7:0];

// Each digit of score
wire [3:0] score_digit0;
wire [3:0] score_digit1;
wire [3:0] score_digit2;
wire [3:0] score_digit3;
wire [3:0] score_digit4;
	
// Update each digit whenever score changes
Score_init(.score(score),.digit4(score_digit4),.digit3(score_digit3),.digit2(score_digit2),.digit1(score_digit1),.digit0(score_digit0));
	
parameter GUI_width = 160; // Width of the GUI
		
// Parameters for weapon
parameter weapon_art_hc = 25; // Horizontal coordinate of Up Left corner of the weapon article
parameter weapon_art_vc = 350; // Vertical coordinate of Up Left corner of the weapon article
parameter weapon_art_width = 108; // Width of weapon article
parameter weapon_art_height = 29; // Height of weapon article

parameter weapon_img0_hc = 63; // Horizontal coordinate of Up Left corner of the weapon image 0
parameter weapon_img0_vc = 416; // Vertical coordinate of Up Left corner of the weapon image 0
parameter weapon_img0_width = 32; // Width of weapon image 0
parameter weapon_img0_height = 32; // Height of weapon image 0

parameter weapon_img1_hc = 55; // Horizontal coordinate of Up Left corner of the weapon image 1
parameter weapon_img1_vc = 408; // Vertical coordinate of Up Left corner of the weapon image 1
parameter weapon_img1_width = 48; // Width of weapon image 1
parameter weapon_img1_height = 48; // Height of weapon image 1

parameter weapon_img2_hc = 48; // Horizontal coordinate of Up Left corner of the weapon image 2
parameter weapon_img2_vc = 400; // Vertical coordinate of Up Left corner of the weapon image 2
parameter weapon_img2_width = 64; // Width of weapon image 2
parameter weapon_img2_height = 64; // Height of weapon image 2

// Curret weapon register
reg[1:0] current_weapon;

		
// Parameters for score		
parameter score_art_hc = 22; // Horizontal coordinate of Up Left corner of the score article
parameter score_art_vc = 69; // Vertical coordinate of Up Left corner of the score article
parameter score_art_width = 115; // Width of score article
parameter score_art_height = 29; // Height of score article
		
parameter score_hc = 19;  // Horizontal coordinate of Up Left corner of the score
parameter score_vc = 109; // Vertical coordinate of Up Left corner of the score
parameter score_width = 24; // Width of each digit of score
parameter score_height = 30; // Height of score
		
// Score register and wires
reg[16:0] score;
	
// Spaceship settings
parameter spaceship_hc = GUI_width + 215;
parameter spaceship_vc = 215;
parameter spaceship_height = 48;
parameter spaceship_width = 48;

wire C_10Hz; 
CLK_10Hz(.CLK(CLK),.CLK_divided(C_10Hz));

// Always block to find the color information of the current location
always @(posedge CLK) begin
	if (~is_blanking & Alive) begin
		pixel = 4'b0000;
		// Check whether we are in the pixels of GUI
		if (hc <= GUI_width) begin 
			if((hc >= score_art_hc) & (vc >= score_art_vc) & (hc <= score_art_hc + score_art_width) & (vc <= score_art_vc + score_art_height)) pixel = GUI_img(hc-score_art_hc,vc-score_art_vc,4'd10);
			else if ((hc >= score_hc) & (vc >= score_vc) & (hc <= score_hc + score_width*5) & (vc <= score_vc + score_height)) begin
				if (hc >= score_hc + 4* score_width) pixel = GUI_img(hc-score_hc-4* score_width,vc-score_vc,score_digit0);
				else if (hc >= score_hc + 3* score_width) pixel = GUI_img(hc-score_hc-3* score_width,vc-score_vc,score_digit1);
				else if (hc >= score_hc + 2* score_width) pixel = GUI_img(hc-score_hc-2* score_width,vc-score_vc,score_digit2);
				else if (hc >= score_hc + score_width) pixel = GUI_img(hc-score_hc- score_width,vc-score_vc,score_digit3);
				else pixel = GUI_img(hc-score_hc-4* score_width,vc-score_vc,score_digit4);
			end
			else if ((hc >= weapon_art_hc) & (vc >= weapon_art_vc) & (hc <= weapon_art_hc + weapon_art_width) & (vc <= weapon_art_vc + weapon_art_height)) pixel = GUI_img(hc-weapon_art_hc,vc-weapon_art_vc,4'd11);
			else if (current_weapon == 2'd0) begin
				if ((hc >= weapon_img0_hc) & (vc >= weapon_img0_vc) & (hc <= weapon_img0_hc + weapon_img0_width) & (vc <= weapon_img0_vc + weapon_img0_height)) pixel = Bullet_img(hc-weapon_img0_hc,vc-weapon_img0_vc,4'd2,2'd0);
			end
			else if (current_weapon == 2'd1) begin
				if ((hc >= weapon_img1_hc) & (vc >= weapon_img1_vc) & (hc <= weapon_img1_hc + weapon_img1_width) & (vc <= weapon_img1_vc + weapon_img1_height)) pixel = Bullet_img(hc-weapon_img1_hc,vc-weapon_img1_vc,4'd2,2'd1);
			end
			else if (current_weapon == 2'd2) begin
				if ((hc >= weapon_img2_hc) & (vc >= weapon_img2_vc) & (hc <= weapon_img2_hc + weapon_img2_width) & (vc <= weapon_img2_vc + weapon_img2_height)) pixel = Bullet_img(hc-weapon_img2_hc,vc-weapon_img2_vc,4'd2,2'd2);
			end
			else pixel = 4'b1111;
		end
		
		else begin
		pixel = pixel_finder();
		end 
	
	end
end

reg is_fire_pressed;
// Unnecessary variable
reg u; 
always @(posedge CLK_10Hz) begin
	if (~RESET) begin
		score = 17'd0;
		Alive = 1'b1;
		enemies_active = 8'd0;
		bullets_active = 32'd0;
	end
	else if (~Fire & ~is_fire_pressed) begin
	is_fire_pressed = 1'b1;
	u = bullet_init(current_weapon,spaceship_angle);
	u = enemies_action();
	u = bullets_action();
	u = enemy_init(rand_mod5_int);
	end
	else if (Alive) begin
	is_fire_pressed = 1'b0;
	u = enemies_action();
	u = bullets_action();
	u = enemy_init(rand_mod5_int);
	end
end


reg [7:0] enemies_dist[7:0];
reg [3:0] enemies_angle[7:0];
reg [3:0] enemies_health[7:0];
reg [3:0] enemies_type[7:0];
reg [7:0]enemies_active;

reg [7:0] bullets_dist[31:0];
reg [3:0] bullets_angle[31:0];
reg [1:0] bullets_type[31:0];
reg [31:0]bullets_active;

reg [3:0] spaceship_angle;

reg temp;

// Always block for updating the state of spaceship
always @(negedge Rotate_CW) spaceship_angle = spaceship_angle + 4'd1;
always @(negedge Rotate_CCW) spaceship_angle = spaceship_angle - 4'd1;

// Always block for updating the type of weapon
always @(negedge Weapon_switch) begin
current_weapon = current_weapon + 2'd1;
if (current_weapon == 2'd3) current_weapon = 2'd0;
end


function [17:0] change_cor(input [7:0] _dist, input [3:0] _angle);
begin
	// cos0 = 1, sin0 = 0
	// cos45 = sin45 = 45/64
	// cos22.5 = 59/64, sin22.5 = 24/64
	// Pozitif y aşağı [17:9]
	// Pozitif x sağ [8:0]
	case(_angle)
		4'd0,4'd4,4'd8,4'd12: begin
			change_cor[8:0] = (_angle == 4'd4) ? 9'd240 -_dist:
				(_angle == 4'd12) ? 9'd240 + _dist
				: 9'd240;
			change_cor[17:9] = (_angle == 4'd0) ? 9'd240 + _dist:
				(_angle == 4'd8) ? 9'd240 - _dist
				: 9'd240;
		end
		4'd2,4'd6,4'd10,4'd14: begin
			reg [14:0] temp1 = 15'd45 * _dist;
			change_cor[8:0] = (_angle == 4'd2 || _angle == 4'd6) ? 9'd240 - temp1[14:6]
			: 9'd240 + temp1[14:6];
			change_cor[17:9] = (_angle == 4'd2 || _angle == 4'd14) ? 9'd240 + temp1[14:6]
			: 9'd240 - temp1[14:6];	
		end
		default: begin
			reg [14:0] temp1 = 15'd59 * _dist;
			reg [14:0] temp2 = 15'd24 * _dist;
			change_cor[8:0] = (_angle == 4'd1 || _angle == 4'd7) ? 9'd240 - temp2[14:6]:
				(_angle == 4'd9 || _angle == 4'd15) ? 9'd240 + temp2[14:6]:
				(_angle == 4'd3 || _angle == 4'd5) ? 9'd240 - temp1[14:6]:
				9'd240 + temp1[14:6];
			change_cor[17:9] = (_angle == 4'd1 || _angle == 4'd15) ? 9'd240 + temp1[14:6]:
				(_angle == 4'd7 || _angle == 4'd9) ? 9'd240 - temp1[14:6]:
				(_angle == 4'd3 || _angle == 4'd13) ? 9'd240 + temp2[14:6]:
				9'd240 - temp2[14:6];
		end
	endcase
end
endfunction

wire[3:0] rand_int;
wire[3:0] rand_mod5_int;

random(CLK_10Hz,rand_int);
random_mod5(CLK_10Hz,rand_mod5_int);

function enemy_init(input [3:0] e_type);
begin
	reg [3:0] i;
	reg stop = 1'b0;
	for(i = 4'd0; i < 4'd8 && ~stop; i = i + 4'd1)
	if(~enemies_active[i]) begin
		stop = 1'b1;
      enemies_active[i] = 1'b1;
		enemies_type[i] = e_type;
		enemies_dist[i] = 8'd240; // Başlangıçta en uzak değer yaptım
		enemies_angle[i] = rand_int; // Random değerini değiştirmek gerek
		enemies_health[i] = (e_type == 0) ? 4'd6:
			(e_type == 1) ? 4'd3:
			(e_type == 2) ? 4'd2:
			(e_type == 3) ? 4'd9:
			4'd15;
	end
end
endfunction


function enemy_move(input [3:0] i);
enemies_dist[i] = (enemies_type[i] == 3'd0) ? enemies_dist[i] - 8'd3 :
	(enemies_type[i] == 3'd1) ? enemies_dist[i] - 8'd4 :
	(enemies_type[i] == 3'd2) ? enemies_dist[i] - 8'd5 :
	(enemies_type[i] == 3'd3) ? enemies_dist[i] - 8'd2 :
	enemies_dist[i] - 8'd1;
endfunction

function enemies_action();
begin
	reg [3:0] i;
	for(i = 4'd0; i < 4'd7; i = i + 4'd1)
	begin
	if (enemies_dist[i] < 5'd24) begin
	enemies_active[i] = 1'b0;
	Alive = 1'b0;
	end
	else if(enemies_active[i]) begin
		temp = enemy_move(i);
	end
	end
end
endfunction

function bullet_init(input [1:0] b_type, input [3:0] angle);
begin
	reg [4:0] i;
	reg [3:0] counter = (b_type == 2'd0) ? 3'd5:
		(b_type == 2'd1) ? 3'd3:
		3'd1;
	
	for(i = 5'd0; i < 5'd31 && counter > 0; i = i + 5'd1)
	if(~bullets_active[i]) begin
        bullets_active[i] = 1'b1;
		bullets_dist[i] = 7'd0; // Başlangıçta merkezde
		bullets_type[i] = b_type;
		bullets_angle[i] = (counter == 5) ? angle + 4'd2:
			(counter == 4) ? angle - 4'd2:
			(counter == 3) ? angle + 4'd1:
			(counter == 2) ? angle - 4'd1:
			angle;
		counter = counter - 1;
	end
end
endfunction

function bullet_move(input [4:0] i);
bullets_dist[i] = (bullets_type[i] == 2'd0) ? bullets_dist[i] + 8'd7 :
	(bullets_type[i] == 2'd1) ? bullets_dist[i] + 8'd5 :
	bullets_dist[i] + 8'd4;
endfunction

function check_col(input [4:0] i);
begin 
	reg [3:0] j;
	reg stop = 1'b0;
	reg [3:0] damage_dealt;
	for(j = 4'd0; j < 4'd7 && ~stop; j = j + 4'd1)
	if(enemies_active[j] && bullets_dist[i] >= enemies_dist[j]) begin
		stop = 1'b1;
		bullets_active[i] = 1'b0; 
		damage_dealt = (bullets_type[i] == 2'd0) ? 4'd2:
			(bullets_type[i] == 2'd1) ? 4'd3: 
			4'd9;
		if(damage_dealt >= enemies_health[j]) begin
			score = (enemies_type[j] == 3'd0) ? score + 17'd6:
				(enemies_type[j] == 3'd1) ? score + 17'd3:
				(enemies_type[j] == 3'd2) ? score + 17'd2:
				(enemies_type[j] == 3'd3) ? score + 17'd9:
				17'd5;
			enemies_active[j] = 1'b0;
		end
		else enemies_health[j] = enemies_health[j] - damage_dealt;
	end
end
endfunction

function bullets_action();
begin
	reg [4:0] i;
	for(i = 5'd0; i < 5'd31; i = i + 5'd1)
	if(bullets_active[i]) begin
		temp = bullet_move(i);
		temp = check_col(i);
	end
end
endfunction

function pixel_finder();
begin
	reg [5:0] i;
	reg [8:0] x;
	reg [8:0] y;
   reg [8:0] d;
	reg [17:0] temp1;
    reg stop = 1'b0;
		
    // For Spaceship
    if(hc >= spaceship_hc && hc <= spaceship_hc + spaceship_width && vc >= spaceship_vc && vc <= spaceship_vc + spaceship_height) begin
		  if (Spaceship_img(hc - spaceship_hc, vc - spaceship_vc, spaceship_angle) != 4'b0000) begin
			  pixel = Spaceship_img(hc - spaceship_hc, vc - spaceship_vc, spaceship_angle);
			  stop = 1'b1;
		  end
    end

	// For enemies
    for (i = 6'd0; i < 6'd7 && ~stop; i = i + 6'd1) begin
			if (enemies_active[i]) begin
			  temp1 = change_cor(enemies_dist[i], enemies_angle[i]);
			  x = temp1[17:9];
			  y = temp1[8:0];

			  d = (enemies_type[i] == 3'd3 | enemies_type[i] == 3'd4) ? 9'd64:
					9'd32;

			  if(hc >= x - d && hc <= x + d && vc >= y - d && vc <= y + d) begin
					if (Enemy_img(hc - x + d, vc - y + d, bullets_angle[i], bullets_type[i]) != 4'b0000) begin
						stop = 1'b1;
						pixel = Enemy_img(hc - x + d, vc - y + d, bullets_angle[i], bullets_type[i]);
					end
			  end
			end
    end

    // For bullets
	for (i = 6'd0; i < 6'd31 && ~stop; i = i + 6'd1) begin
		if (bullets_active[i]) begin
			  temp1 = change_cor(bullets_dist[i], bullets_angle[i]);
			  x = temp1[17:9] + GUI_width;
			  y = temp1[8:0];

			  d = (bullets_type[i] == 3'd0) ? 9'd16:
					(bullets_type[i] == 3'd1) ? 9'd24:
					9'd32; 

			  if(hc >= x - d && hc <= x + d && vc >= y - d && vc <= y + d) begin
					if(Bullet_img(hc - x + d, vc - y + d, bullets_angle[i], bullets_type[i]) != 4'b0000) begin
						stop = 1'b1;
						pixel = Bullet_img(hc - x + d, vc - y + d, bullets_angle[i], bullets_type[i]);
					end
			  end
		end
    end
end
endfunction

function [3:0] Spaceship_img(input [6:0] x, input [6:0] y, input [3:0] angle);
begin
//case(angle)
//// Spaceship 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//endcase
//end
//// Spaceship 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10,6'd13,6'd14: Spaceship_img = 4'd13;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Spaceship_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd10,6'd13,6'd14,6'd15: Spaceship_img = 4'd13;
//6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25: Spaceship_img = 4'd3;
//6'd13,6'd14,6'd15,6'd17,6'd18,6'd19: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd16: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd3;
//6'd45: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd22,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd14;
//6'd39: Spaceship_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd3;
//6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24: Spaceship_img = 4'd3;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd14;
//6'd27: Spaceship_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd28,6'd29,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd30,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//6'd1,6'd2,6'd3,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//6'd1,6'd6,6'd7,6'd8,6'd9,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd32: Spaceship_img = 4'd13;
//6'd16,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd10,6'd26,6'd41,6'd42: Spaceship_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd4,6'd8,6'd9,6'd10,6'd24,6'd25,6'd26,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd12,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd5,6'd6,6'd7: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd3,6'd4,6'd5,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd8,6'd11: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd10;
//6'd22,6'd23,6'd24,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd9,6'd10,6'd11,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd13,6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd27,6'd28,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd26,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd10,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd33: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd17,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd33,6'd34: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd13,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd15,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30: Spaceship_img = 4'd3;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd28: Spaceship_img = 4'd13;
//6'd12,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd11,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd3;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd12;
//6'd9,6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd12;
//6'd10,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd12;
//6'd9,6'd10,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd23: Spaceship_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//endcase
//end
//// Spaceship 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd14,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd13;
//6'd18,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd24,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd23,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd14: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd16,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd12: Spaceship_img = 4'd2;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd16,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13: Spaceship_img = 4'd2;
//6'd14: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd14,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd15,6'd20,6'd21,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//6'd33: Spaceship_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd38,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd35: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd44,6'd45,6'd46,6'd47: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd13: Spaceship_img = 4'd2;
//6'd14: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd43,6'd44,6'd47,6'd48: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11: Spaceship_img = 4'd0;
//6'd12: Spaceship_img = 4'd2;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13: Spaceship_img = 4'd0;
//6'd14: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd27,6'd28,6'd29,6'd30,6'd35,6'd39: Spaceship_img = 4'd13;
//6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd43,6'd44,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd22,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd46: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd29: Spaceship_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20: Spaceship_img = 4'd10;
//6'd16,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd18,6'd22,6'd23,6'd24,6'd25,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd18,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd14,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd31,6'd35,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd33,6'd37: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd24,6'd25: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd29,6'd33: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd13,6'd14,6'd24,6'd25,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd31,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd24,6'd25,6'd32,6'd33,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd37,6'd38: Spaceship_img = 4'd3;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd3;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Spaceship_img = 4'd13;
//6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd30,6'd36: Spaceship_img = 4'd2;
//6'd28,6'd29,6'd37,6'd38: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd41,6'd42,6'd45,6'd46: Spaceship_img = 4'd13;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd37: Spaceship_img = 4'd2;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd13;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd12;
//6'd16: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd12;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10: Spaceship_img = 4'd12;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//endcase
//end
//// Spaceship 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd23: Spaceship_img = 4'd14;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd6,6'd7,6'd22,6'd23,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd22,6'd23,6'd24,6'd41,6'd44,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd21,6'd22,6'd23,6'd24,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd12,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd23,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd24,6'd25,6'd26,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd40,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd24,6'd25,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd26,6'd33,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd31,6'd32,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd23,6'd24,6'd25,6'd36,6'd37: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd32,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd38,6'd39,6'd40,6'd43,6'd44: Spaceship_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd17,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd24,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd18,6'd27,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd19,6'd39,6'd40,6'd41: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd13: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd44,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11: Spaceship_img = 4'd0;
//6'd12,6'd13,6'd14: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd13,6'd14: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd0;
//6'd21,6'd22: Spaceship_img = 4'd10;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd39,6'd46: Spaceship_img = 4'd14;
//6'd15: Spaceship_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40: Spaceship_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd10;
//6'd17,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd26,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39,6'd40,6'd41: Spaceship_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd10;
//6'd17,6'd18,6'd19,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd44,6'd45: Spaceship_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39,6'd40,6'd41: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38: Spaceship_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd41: Spaceship_img = 4'd3;
//6'd25: Spaceship_img = 4'd10;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd16,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd33,6'd34: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd33: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd24: Spaceship_img = 4'd13;
//6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd23,6'd24,6'd25: Spaceship_img = 4'd13;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd23,6'd24,6'd25: Spaceship_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd13: Spaceship_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd12;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd12;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18: Spaceship_img = 4'd12;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//endcase
//end
//// Spaceship 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//6'd1,6'd2,6'd3,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//6'd1,6'd2,6'd3,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//6'd1,6'd2,6'd3,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd40,6'd41,6'd42: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd40,6'd41,6'd42: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd40,6'd41,6'd42: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//endcase
//end
//// Spaceship 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd26,6'd27,6'd42,6'd43: Spaceship_img = 4'd13;
//6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd5,6'd8,6'd25,6'd26,6'd27,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd13;
//6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd25,6'd26,6'd27,6'd28,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd3,6'd4,6'd5,6'd6,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd26,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd23,6'd24,6'd25,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd9,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd24,6'd25,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd16,6'd23,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd22,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd17,6'd18,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd24,6'd25,6'd26,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd13,6'd14,6'd17,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd3;
//6'd5,6'd6,6'd9,6'd10,6'd11,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd32,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd17,6'd18,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd16,6'd25,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd22,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd10,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd8,6'd9,6'd10,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd36: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd13,6'd14: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd5,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd37: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd35,6'd36: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28: Spaceship_img = 4'd10;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd3,6'd10,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//6'd34: Spaceship_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9: Spaceship_img = 4'd3;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//6'd20,6'd21,6'd22,6'd32: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd23,6'd30,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10: Spaceship_img = 4'd3;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//6'd20,6'd21,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10: Spaceship_img = 4'd3;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd10;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd11,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd17: Spaceship_img = 4'd3;
//6'd24: Spaceship_img = 4'd10;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd19,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd25,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd36: Spaceship_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//6'd26: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32: Spaceship_img = 4'd12;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//endcase
//end
//// Spaceship 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd18,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd18,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd18,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd20,6'd25,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd26,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd18,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd37: Spaceship_img = 4'd2;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd20,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd36: Spaceship_img = 4'd2;
//6'd35: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd28,6'd29,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd14;
//6'd16: Spaceship_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd11,6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//6'd14,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd4,6'd5,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd36: Spaceship_img = 4'd2;
//6'd35: Spaceship_img = 4'd3;
//6'd1,6'd2,6'd5,6'd6,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd11,6'd12,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd37: Spaceship_img = 4'd2;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd9,6'd10,6'd11,6'd13,6'd14,6'd15,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd35: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd10,6'd14,6'd19,6'd20,6'd21,6'd22,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd5,6'd6,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd27,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd3,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29: Spaceship_img = 4'd10;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd33: Spaceship_img = 4'd12;
//6'd8,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd9,6'd24,6'd25,6'd26,6'd27,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd11,6'd12,6'd13,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21,6'd22,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd35: Spaceship_img = 4'd13;
//6'd10,6'd14,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//6'd12,6'd16,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd9,6'd10,6'd11,6'd13,6'd14,6'd15,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd10;
//6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd16,6'd20,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27: Spaceship_img = 4'd10;
//6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd19,6'd20,6'd21,6'd24,6'd25,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd3,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd16,6'd17,6'd24,6'd25,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd15: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd14: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd19: Spaceship_img = 4'd2;
//6'd11,6'd12,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd7,6'd8,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd12,6'd20: Spaceship_img = 4'd2;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Spaceship_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd12;
//6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Spaceship_img = 4'd12;
//6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39: Spaceship_img = 4'd12;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//endcase
//end
//// Spaceship 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd12;
//6'd9,6'd10,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd23: Spaceship_img = 4'd14;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd12;
//6'd10,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd3;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd12;
//6'd9,6'd10,6'd11,6'd12,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd3;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd11,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30: Spaceship_img = 4'd3;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd28: Spaceship_img = 4'd13;
//6'd12,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd15,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd13,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd33,6'd34: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd33: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd17,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd27,6'd28,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd26,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd10,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd13,6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd10;
//6'd22,6'd23,6'd24,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd9,6'd10,6'd11,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd3,6'd4,6'd5,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd8,6'd11: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd12,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd5,6'd6,6'd7: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd4,6'd8,6'd9,6'd10,6'd24,6'd25,6'd26,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd10,6'd26,6'd41,6'd42: Spaceship_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd6,6'd7,6'd8,6'd9,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd32: Spaceship_img = 4'd13;
//6'd16,6'd19,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd2,6'd3,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd20,6'd21: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd28,6'd29,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd30,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24: Spaceship_img = 4'd3;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd14;
//6'd27: Spaceship_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd3;
//6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd3;
//6'd45: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd22,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd14;
//6'd39: Spaceship_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25: Spaceship_img = 4'd3;
//6'd13,6'd14,6'd15,6'd17,6'd18,6'd19: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd16: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd10,6'd13,6'd14,6'd15: Spaceship_img = 4'd13;
//6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Spaceship_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10,6'd13,6'd14: Spaceship_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//endcase
//end
//// Spaceship 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39: Spaceship_img = 4'd12;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Spaceship_img = 4'd12;
//6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd12;
//6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd12,6'd20: Spaceship_img = 4'd2;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Spaceship_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd19: Spaceship_img = 4'd2;
//6'd11,6'd12,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd7,6'd8,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd14: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//6'd1,6'd2,6'd16,6'd17,6'd24,6'd25,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd15: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//6'd1,6'd2,6'd3,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd11,6'd12: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27: Spaceship_img = 4'd10;
//6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd19,6'd20,6'd21,6'd24,6'd25,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd10;
//6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd16,6'd20,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//6'd12,6'd16,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd9,6'd10,6'd11,6'd13,6'd14,6'd15,6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd11,6'd12,6'd13,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21,6'd22,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd35: Spaceship_img = 4'd13;
//6'd10,6'd14,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd10;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd9,6'd24,6'd25,6'd26,6'd27,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29: Spaceship_img = 4'd10;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd33: Spaceship_img = 4'd12;
//6'd8,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd3,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd5,6'd6,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd27,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd35: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd10,6'd14,6'd19,6'd20,6'd21,6'd22,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd9,6'd10,6'd11,6'd13,6'd14,6'd15,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd37: Spaceship_img = 4'd2;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd36: Spaceship_img = 4'd2;
//6'd35: Spaceship_img = 4'd3;
//6'd1,6'd2,6'd5,6'd6,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd11,6'd12,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//6'd14,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd2,6'd3,6'd4,6'd5,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd11,6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd14;
//6'd16: Spaceship_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd28,6'd29,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd36: Spaceship_img = 4'd2;
//6'd35: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd37: Spaceship_img = 4'd2;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd20,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd18,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd26,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd20,6'd25,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd18,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd18,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd18,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd18: Spaceship_img = 4'd14;
//endcase
//end
//endcase
//end
//// Spaceship 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32: Spaceship_img = 4'd12;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd12;
//6'd26: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd36: Spaceship_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd25,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd19,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd17: Spaceship_img = 4'd3;
//6'd24: Spaceship_img = 4'd10;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10: Spaceship_img = 4'd3;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd10;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd11,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10: Spaceship_img = 4'd3;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//6'd20,6'd21,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9: Spaceship_img = 4'd3;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd10;
//6'd20,6'd21,6'd22,6'd32: Spaceship_img = 4'd12;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd23,6'd30,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd27,6'd28: Spaceship_img = 4'd10;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd3,6'd10,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//6'd34: Spaceship_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd35,6'd36: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd37: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd5,6'd26,6'd27,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd36: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd13,6'd14: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd8,6'd9,6'd10,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd10,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd22,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd17,6'd18,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd16,6'd25,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd32,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38,6'd39,6'd40: Spaceship_img = 4'd3;
//6'd5,6'd6,6'd9,6'd10,6'd11,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd13,6'd14,6'd17,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd17,6'd18,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd24,6'd25,6'd26,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd22,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd4,6'd5,6'd6,6'd9,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd24,6'd25,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd16,6'd23,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd3,6'd4,6'd5,6'd6,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd26,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd23,6'd24,6'd25,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd25,6'd26,6'd27,6'd28,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd5,6'd8,6'd25,6'd26,6'd27,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd13;
//6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd3,6'd4,6'd26,6'd27,6'd42,6'd43: Spaceship_img = 4'd13;
//6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd26,6'd27: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//endcase
//end
//// Spaceship 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd40,6'd41,6'd42: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd40,6'd41,6'd42: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd40,6'd41,6'd42: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd3,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10,6'd11,6'd12,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//endcase
//end
//endcase
//end
//// Spaceship 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18: Spaceship_img = 4'd12;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd12;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd12;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//6'd13: Spaceship_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd23,6'd24,6'd25: Spaceship_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd23,6'd24,6'd25: Spaceship_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd33: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd24: Spaceship_img = 4'd13;
//6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd33,6'd34: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd32,6'd41: Spaceship_img = 4'd3;
//6'd25: Spaceship_img = 4'd10;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//6'd16,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34: Spaceship_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39,6'd40,6'd41: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38: Spaceship_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39,6'd40,6'd41: Spaceship_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd10;
//6'd17,6'd18,6'd19,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd44,6'd45: Spaceship_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40: Spaceship_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Spaceship_img = 4'd10;
//6'd17,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd26,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd0;
//6'd21,6'd22: Spaceship_img = 4'd10;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd39,6'd46: Spaceship_img = 4'd14;
//6'd15: Spaceship_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd13,6'd14: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11: Spaceship_img = 4'd0;
//6'd12,6'd13,6'd14: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd44,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd13: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd27,6'd28: Spaceship_img = 4'd13;
//6'd19,6'd39,6'd40,6'd41: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd18,6'd27,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd24,6'd33: Spaceship_img = 4'd13;
//6'd17,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd15,6'd16,6'd17,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd38,6'd39,6'd40,6'd43,6'd44: Spaceship_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd25,6'd32,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd31,6'd32,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd23,6'd24,6'd25,6'd36,6'd37: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd40,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd24,6'd25,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd26,6'd33,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd12;
//6'd8,6'd9,6'd10,6'd23,6'd40,6'd41,6'd42: Spaceship_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd24,6'd25,6'd26,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd21,6'd22,6'd23,6'd24,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd12,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd22,6'd23,6'd24,6'd41,6'd44,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd6,6'd7,6'd22,6'd23,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//6'd23: Spaceship_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd12;
//endcase
//end
//endcase
//end
//// Spaceship 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd10: Spaceship_img = 4'd12;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd9,6'd10,6'd11: Spaceship_img = 4'd12;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd12;
//6'd16: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19: Spaceship_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd29,6'd37: Spaceship_img = 4'd2;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd30,6'd36: Spaceship_img = 4'd2;
//6'd28,6'd29,6'd37,6'd38: Spaceship_img = 4'd3;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd41,6'd42,6'd45,6'd46: Spaceship_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd3;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Spaceship_img = 4'd13;
//6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd24,6'd25,6'd32,6'd33,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd37,6'd38: Spaceship_img = 4'd3;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd13,6'd14,6'd24,6'd25,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd31,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd29,6'd33: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd33,6'd37: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd24,6'd25: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd18,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd14,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd13;
//6'd31,6'd35,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Spaceship_img = 4'd12;
//6'd18,6'd22,6'd23,6'd24,6'd25,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20: Spaceship_img = 4'd10;
//6'd16,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd46: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd29: Spaceship_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd43,6'd44,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd22,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13: Spaceship_img = 4'd0;
//6'd14: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd27,6'd28,6'd29,6'd30,6'd35,6'd39: Spaceship_img = 4'd13;
//6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//default: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11: Spaceship_img = 4'd0;
//6'd12: Spaceship_img = 4'd2;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Spaceship_img = 4'd0;
//6'd13: Spaceship_img = 4'd2;
//6'd14: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd43,6'd44,6'd47,6'd48: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd35: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd44,6'd45,6'd46,6'd47: Spaceship_img = 4'd13;
//default: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd45,6'd46: Spaceship_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd38,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd20: Spaceship_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//6'd33: Spaceship_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd15,6'd20,6'd21,6'd30,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd14,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13: Spaceship_img = 4'd2;
//6'd14: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd12: Spaceship_img = 4'd2;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd16,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd13,6'd14,6'd15: Spaceship_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd16,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd14: Spaceship_img = 4'd3;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd23,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd24,6'd29: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16: Spaceship_img = 4'd13;
//6'd17,6'd18,6'd19,6'd30,6'd31,6'd32: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17: Spaceship_img = 4'd13;
//6'd18,6'd31: Spaceship_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd16,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd15,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd14,6'd31: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd31: Spaceship_img = 4'd14;
//endcase
//end
//endcase
//end
//// Spaceship 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd34,6'd35,6'd36,6'd39: Spaceship_img = 4'd13;
//6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25: Spaceship_img = 4'd3;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd33,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd3;
//6'd4: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd27,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//6'd10: Spaceship_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd3;
//6'd4,6'd5,6'd6: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25: Spaceship_img = 4'd3;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//6'd22: Spaceship_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd1,6'd2,6'd20,6'd21,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd19: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//6'd1,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd30: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//6'd1,6'd40,6'd41,6'd42,6'd43,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd17,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//6'd1,6'd2,6'd3: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5: Spaceship_img = 4'd0;
//6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd23,6'd39,6'd46,6'd47: Spaceship_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd48: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd23,6'd24,6'd25,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47: Spaceship_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd42,6'd43,6'd44: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd44,6'd45,6'd46,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd38,6'd41,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd13,6'd14,6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd38,6'd39,6'd40,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd36: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd21,6'd22,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd23,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd15,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd32: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd24,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd34: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20: Spaceship_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd21: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd38: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd3;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd39: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd39,6'd40: Spaceship_img = 4'd13;
//6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//endcase
//end
//// Spaceship 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27,6'd40,6'd41,6'd42: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd43,6'd44,6'd45: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Spaceship_img = 4'd12;
//6'd25,6'd26,6'd27,6'd46,6'd47,6'd48: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd3;
//6'd28,6'd29,6'd30: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//endcase
//end
//endcase
//end
//// Spaceship 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd1: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd38: Spaceship_img = 4'd12;
//6'd23,6'd24,6'd25,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//6'd22: Spaceship_img = 4'd14;
//endcase
//end
//6'd3: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd39,6'd40: Spaceship_img = 4'd13;
//6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd5: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd39: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd37,6'd38,6'd39: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26: Spaceship_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20: Spaceship_img = 4'd3;
//6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23,6'd24,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd12;
//6'd22,6'd23,6'd38: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd19,6'd20: Spaceship_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Spaceship_img = 4'd12;
//6'd21: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd34: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd20,6'd21,6'd22,6'd33,6'd34,6'd35: Spaceship_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd24,6'd25,6'd26,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd17: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd24,6'd34,6'd35,6'd36: Spaceship_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd31,6'd32,6'd33: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd19,6'd20,6'd21,6'd32,6'd33,6'd34: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24: Spaceship_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16: Spaceship_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd32: Spaceship_img = 4'd13;
//6'd22,6'd23,6'd24,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Spaceship_img = 4'd12;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd17,6'd18,6'd19,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Spaceship_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd16,6'd17,6'd21,6'd22,6'd24,6'd25,6'd26: Spaceship_img = 4'd12;
//6'd18,6'd19,6'd20,6'd23,6'd27,6'd28,6'd29: Spaceship_img = 4'd13;
//6'd15,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd15,6'd16,6'd17,6'd24,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd13,6'd14,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd36: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd15,6'd16,6'd17,6'd25,6'd26,6'd27: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd13,6'd14,6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd13;
//6'd31,6'd32,6'd33,6'd38,6'd39,6'd40,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd44,6'd45,6'd46,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd16,6'd17,6'd18,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd38,6'd41,6'd42,6'd43: Spaceship_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd48: Spaceship_img = 4'd0;
//6'd19,6'd20,6'd21: Spaceship_img = 4'd10;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd42,6'd43,6'd44: Spaceship_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd48: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd9,6'd10,6'd23,6'd24,6'd25,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47: Spaceship_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6: Spaceship_img = 4'd0;
//6'd20,6'd21,6'd22: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd7,6'd8,6'd23,6'd39,6'd46,6'd47: Spaceship_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5: Spaceship_img = 4'd0;
//6'd20,6'd21: Spaceship_img = 4'd10;
//default: Spaceship_img = 4'd12;
//6'd22,6'd23: Spaceship_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd21,6'd22,6'd23: Spaceship_img = 4'd13;
//6'd27,6'd28,6'd29: Spaceship_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd40,6'd41,6'd42,6'd43,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd17,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd30,6'd33: Spaceship_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//default: Spaceship_img = 4'd12;
//6'd15,6'd16,6'd17,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd30: Spaceship_img = 4'd13;
//6'd28,6'd29,6'd31,6'd32,6'd33,6'd34: Spaceship_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd20,6'd21,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Spaceship_img = 4'd0;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd19: Spaceship_img = 4'd12;
//default: Spaceship_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Spaceship_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd25: Spaceship_img = 4'd3;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Spaceship_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//6'd22: Spaceship_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25: Spaceship_img = 4'd3;
//6'd4,6'd5,6'd6: Spaceship_img = 4'd12;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Spaceship_img = 4'd3;
//6'd4: Spaceship_img = 4'd12;
//6'd11,6'd12,6'd27,6'd30,6'd31,6'd32: Spaceship_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Spaceship_img = 4'd14;
//6'd10: Spaceship_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd24,6'd25: Spaceship_img = 4'd3;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36: Spaceship_img = 4'd13;
//6'd33,6'd37,6'd38,6'd39: Spaceship_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd34,6'd35,6'd36,6'd39: Spaceship_img = 4'd13;
//6'd37,6'd38: Spaceship_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd31,6'd32,6'd33: Spaceship_img = 4'd3;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Spaceship_img = 4'd13;
//endcase
//end
//6'd41: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd35,6'd36,6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39,6'd40,6'd41: Spaceship_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Spaceship_img = 4'd0;
//6'd39: Spaceship_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Spaceship_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase


end
endfunction



function [3:0] Enemy_img(input [6:0] x, input [6:0] y, input [3:0] angle, input [2:0] e_type);
begin

//case(e_type)
//
//2'd0: begin
//case(angle)
//// Enemy_type_0 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd13;
//6'd22,6'd23,6'd25,6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd25,6'd26,6'd27: Enemy_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd13;
//6'd21,6'd22,6'd26,6'd27: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd13;
//6'd21,6'd22,6'd26,6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd4;
//6'd21,6'd22,6'd23,6'd24: Enemy_img = 4'd13;
//6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd4;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd20,6'd21: Enemy_img = 4'd4;
//6'd18,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17,6'd18: Enemy_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd27,6'd31: Enemy_img = 4'd9;
//6'd45: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd25,6'd29,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd26,6'd30: Enemy_img = 4'd9;
//6'd19,6'd20,6'd24,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd26,6'd30: Enemy_img = 4'd10;
//6'd18,6'd19,6'd20,6'd24,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd26,6'd30: Enemy_img = 4'd9;
//6'd18,6'd19,6'd20,6'd24,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd26,6'd30: Enemy_img = 4'd9;
//6'd19,6'd20,6'd24,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd20,6'd21,6'd25,6'd29,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd45: Enemy_img = 4'd14;
//6'd18,6'd23,6'd27,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd16,6'd17,6'd24,6'd25,6'd26,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17,6'd18: Enemy_img = 4'd3;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd20,6'd21: Enemy_img = 4'd3;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd18,6'd22,6'd29,6'd33,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd3;
//6'd19,6'd20,6'd21,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd18,6'd26,6'd27,6'd28,6'd29,6'd33,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd31,6'd32,6'd37,6'd38: Enemy_img = 4'd14;
//6'd19,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd19: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd19,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//6'd20,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Enemy_img = 4'd14;
//6'd20,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Enemy_img = 4'd14;
//6'd20,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd14;
//6'd21,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd14;
//6'd21,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd14;
//6'd21,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//6'd22,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//6'd22,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//6'd23,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//6'd23,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16: Enemy_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16: Enemy_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16,6'd17,6'd18: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd18: Enemy_img = 4'd13;
//6'd16,6'd17,6'd19,6'd20,6'd21: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd18: Enemy_img = 4'd13;
//6'd16,6'd17,6'd19,6'd20,6'd21,6'd22,6'd23,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd3;
//6'd18,6'd19,6'd20: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd3;
//6'd18,6'd19,6'd20,6'd21: Enemy_img = 4'd13;
//6'd16,6'd17,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd29,6'd30,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Enemy_img = 4'd13;
//6'd16,6'd17,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd43,6'd47: Enemy_img = 4'd13;
//6'd16,6'd17,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd44,6'd45,6'd46: Enemy_img = 4'd13;
//6'd16,6'd17,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd4;
//6'd19,6'd20,6'd21,6'd42,6'd43,6'd44: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd4;
//6'd19,6'd20,6'd40,6'd41: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd21,6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23: Enemy_img = 4'd4;
//6'd18,6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd16,6'd17,6'd19,6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd9;
//6'd35,6'd36: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19: Enemy_img = 4'd4;
//6'd32,6'd33,6'd34: Enemy_img = 4'd13;
//6'd17,6'd18,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd31,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17,6'd18: Enemy_img = 4'd4;
//6'd26,6'd29: Enemy_img = 4'd9;
//6'd31,6'd32: Enemy_img = 4'd13;
//6'd16,6'd19,6'd20,6'd21,6'd23,6'd24,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd41,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17: Enemy_img = 4'd3;
//6'd22,6'd25,6'd30: Enemy_img = 4'd9;
//6'd28: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd24,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16: Enemy_img = 4'd3;
//6'd22,6'd30: Enemy_img = 4'd9;
//6'd26: Enemy_img = 4'd10;
//6'd17,6'd18,6'd19,6'd20,6'd24,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd26: Enemy_img = 4'd9;
//6'd24: Enemy_img = 4'd13;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd28,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd32,6'd39,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd9;
//6'd22: Enemy_img = 4'd10;
//6'd20: Enemy_img = 4'd13;
//6'd19,6'd24,6'd30,6'd31,6'd35,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd28,6'd33,6'd34,6'd39,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd9;
//6'd18,6'd19: Enemy_img = 4'd13;
//6'd20,6'd21,6'd25,6'd26,6'd29,6'd30,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd31,6'd32,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd3;
//6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd24,6'd26,6'd27,6'd31,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd26,6'd31,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd3;
//6'd21,6'd22,6'd23,6'd26,6'd27,6'd28: Enemy_img = 4'd14;
//6'd20,6'd24,6'd25,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd3;
//6'd20,6'd21,6'd22,6'd23,6'd25,6'd32,6'd33: Enemy_img = 4'd14;
//6'd19,6'd24,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26: Enemy_img = 4'd3;
//6'd24,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd18,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd21,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd21,6'd22,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd23,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd23,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd25,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd27,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd14;
//6'd29,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd14;
//6'd30,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//6'd25,6'd26,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd26,6'd32,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd26,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36: Enemy_img = 4'd14;
//6'd27,6'd35,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd27,6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42: Enemy_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd28,6'd40,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd41: Enemy_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd3;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd39,6'd40,6'd41,6'd42,6'd44: Enemy_img = 4'd14;
//6'd28,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd35: Enemy_img = 4'd3;
//6'd45: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd34,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd28,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd3;
//6'd44: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd35,6'd36,6'd42,6'd43,6'd46,6'd48: Enemy_img = 4'd14;
//6'd28,6'd34,6'd37,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd48: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd9;
//6'd43: Enemy_img = 4'd13;
//6'd29,6'd30,6'd34,6'd35,6'd36,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd28,6'd33,6'd37,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd47,6'd48: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd10;
//6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd28,6'd32,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd40,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd33,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd47: Enemy_img = 4'd4;
//6'd38,6'd42,6'd43: Enemy_img = 4'd9;
//6'd30,6'd31,6'd34,6'd41,6'd44,6'd45,6'd46,6'd48: Enemy_img = 4'd14;
//6'd28,6'd29,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd46: Enemy_img = 4'd4;
//6'd39: Enemy_img = 4'd10;
//6'd33,6'd35,6'd36,6'd37,6'd41,6'd44,6'd45,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd46: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd9;
//6'd38: Enemy_img = 4'd13;
//6'd28,6'd29,6'd32,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd26,6'd27,6'd30,6'd31,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd45: Enemy_img = 4'd4;
//6'd35,6'd36,6'd40: Enemy_img = 4'd9;
//6'd48: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd38,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd9;
//6'd36: Enemy_img = 4'd10;
//6'd47,6'd48: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd23,6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd9;
//6'd34,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd45,6'd50,6'd51: Enemy_img = 4'd14;
//6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43: Enemy_img = 4'd4;
//6'd33,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd51,6'd52: Enemy_img = 4'd14;
//6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42: Enemy_img = 4'd4;
//6'd32,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd43,6'd52,6'd53: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd4;
//6'd31,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd45,6'd52,6'd53: Enemy_img = 4'd14;
//6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd4;
//6'd30,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd4;
//6'd29,6'd52: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54: Enemy_img = 4'd14;
//6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd27: Enemy_img = 4'd13;
//6'd25,6'd26,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd26: Enemy_img = 4'd13;
//6'd24,6'd25,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd53,6'd55: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd25,6'd27: Enemy_img = 4'd13;
//6'd23,6'd24,6'd29,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd27: Enemy_img = 4'd13;
//6'd22,6'd23,6'd28,6'd33,6'd34: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd13;
//6'd22,6'd32,6'd33: Enemy_img = 4'd14;
//6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd36: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd3;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd39,6'd44: Enemy_img = 4'd14;
//6'd19,6'd20,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd44: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd43: Enemy_img = 4'd14;
//6'd20: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd44: Enemy_img = 4'd3;
//6'd39,6'd40: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd21,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd3;
//6'd44: Enemy_img = 4'd4;
//6'd39: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd35,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46: Enemy_img = 4'd14;
//6'd22,6'd23,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd3;
//6'd44: Enemy_img = 4'd4;
//6'd36,6'd37,6'd38: Enemy_img = 4'd9;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd41,6'd42,6'd43,6'd45,6'd46: Enemy_img = 4'd14;
//6'd33,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd3;
//6'd44: Enemy_img = 4'd4;
//6'd39: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd33,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd23,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd9;
//6'd38,6'd46: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd31,6'd32,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48: Enemy_img = 4'd14;
//6'd24,6'd25,6'd30,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd44: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd9;
//6'd46: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd31,6'd32,6'd39,6'd42,6'd43,6'd45,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd24,6'd30,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd43,6'd44: Enemy_img = 4'd4;
//6'd36: Enemy_img = 4'd9;
//6'd37: Enemy_img = 4'd10;
//6'd46,6'd47,6'd48: Enemy_img = 4'd13;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd39,6'd40,6'd41,6'd42,6'd45,6'd49,6'd50: Enemy_img = 4'd14;
//6'd25,6'd29,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd38: Enemy_img = 4'd9;
//6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd29,6'd32,6'd34,6'd40,6'd41,6'd42,6'd44,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd14;
//6'd25,6'd26,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd38: Enemy_img = 4'd9;
//6'd36,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd35,6'd37,6'd40,6'd41,6'd42,6'd44,6'd45,6'd51,6'd52,6'd53: Enemy_img = 4'd14;
//6'd25,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd34: Enemy_img = 4'd9;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd39,6'd40,6'd41,6'd42,6'd44,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd36: Enemy_img = 4'd9;
//6'd35: Enemy_img = 4'd10;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd13;
//6'd31,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd42,6'd43: Enemy_img = 4'd4;
//6'd45,6'd46,6'd47,6'd48,6'd50: Enemy_img = 4'd13;
//6'd27,6'd28,6'd31,6'd33,6'd34,6'd38,6'd39,6'd40,6'd41,6'd44,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd26,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd9;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd34: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd53,6'd55: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd34: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42: Enemy_img = 4'd4;
//6'd33: Enemy_img = 4'd13;
//6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44: Enemy_img = 4'd14;
//6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42: Enemy_img = 4'd4;
//6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd24,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd4;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd24,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd32: Enemy_img = 4'd13;
//6'd25,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd32: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd31: Enemy_img = 4'd13;
//6'd29,6'd30,6'd32,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd13;
//6'd29,6'd30,6'd32,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd28,6'd29,6'd31,6'd32,6'd37,6'd38: Enemy_img = 4'd14;
//6'd25,6'd26,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd27,6'd29,6'd31,6'd33,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd28,6'd29,6'd33,6'd37: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd13;
//6'd28,6'd32: Enemy_img = 4'd14;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd13;
//6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd13;
//6'd27: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd39: Enemy_img = 4'd3;
//6'd38: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd39: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd31,6'd34,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//6'd28,6'd29,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd4;
//6'd43: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd37,6'd38,6'd39,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd19,6'd20,6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd4;
//6'd33,6'd34,6'd36: Enemy_img = 4'd9;
//6'd35: Enemy_img = 4'd10;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd38,6'd39,6'd40,6'd42,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd17,6'd18,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd9;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd39,6'd40,6'd42,6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd15,6'd16,6'd30,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd32,6'd37,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd4;
//6'd35,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//default: Enemy_img = 4'd14;
//6'd13,6'd14,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd4;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd32,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd15,6'd16,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd33,6'd34,6'd36: Enemy_img = 4'd9;
//6'd35: Enemy_img = 4'd10;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd38,6'd39,6'd40,6'd41,6'd43,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd17,6'd18,6'd28,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd9;
//6'd44,6'd45,6'd46: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd39,6'd40,6'd41,6'd43,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd19,6'd20,6'd28,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd35,6'd44: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd33,6'd34,6'd36,6'd38,6'd39,6'd40,6'd41,6'd43,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd21,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd24,6'd25,6'd26,6'd31,6'd32,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd22,6'd23,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd33,6'd34,6'd36: Enemy_img = 4'd9;
//6'd35: Enemy_img = 4'd10;
//6'd25,6'd26,6'd28,6'd29,6'd31,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd23,6'd24,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd9;
//6'd27,6'd28,6'd29,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd24,6'd25,6'd30,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd31,6'd33,6'd34,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44: Enemy_img = 4'd14;
//6'd25,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd43: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd43: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd43: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd43: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd33,6'd34,6'd36,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd33,6'd34,6'd36,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27,6'd31,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd33,6'd34,6'd36,6'd42: Enemy_img = 4'd14;
//6'd27,6'd31,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd33,6'd34,6'd36,6'd38: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd33,6'd34,6'd36,6'd38: Enemy_img = 4'd14;
//6'd30,6'd31,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd37: Enemy_img = 4'd13;
//6'd32,6'd34,6'd38: Enemy_img = 4'd14;
//6'd30,6'd31,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd3;
//6'd31,6'd34,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd3;
//6'd34: Enemy_img = 4'd4;
//6'd32,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd4;
//6'd29,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd39,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd4;
//6'd29,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd13;
//6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd4;
//6'd30,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd36,6'd37: Enemy_img = 4'd4;
//6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd33,6'd34,6'd35,6'd38,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd37: Enemy_img = 4'd4;
//6'd31,6'd32,6'd33: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd40,6'd41,6'd42: Enemy_img = 4'd13;
//6'd23,6'd25,6'd26,6'd27,6'd35,6'd36,6'd38,6'd39,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd37,6'd38: Enemy_img = 4'd4;
//6'd29: Enemy_img = 4'd9;
//6'd41,6'd42: Enemy_img = 4'd13;
//6'd22,6'd23,6'd25,6'd26,6'd27,6'd34,6'd35,6'd36,6'd39,6'd40,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd20,6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd4;
//6'd31,6'd41: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd25,6'd26,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd39: Enemy_img = 4'd4;
//6'd33: Enemy_img = 4'd9;
//6'd20,6'd21,6'd22,6'd23,6'd25,6'd29,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd18,6'd19,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd4;
//6'd31,6'd34: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26,6'd29,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd27,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd40,6'd41: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd9;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd34,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43: Enemy_img = 4'd14;
//6'd15,6'd16,6'd17,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd33: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd31,6'd32,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43: Enemy_img = 4'd14;
//6'd15,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd34: Enemy_img = 4'd9;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd14,6'd15,6'd26,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd42: Enemy_img = 4'd4;
//6'd32,6'd33,6'd36: Enemy_img = 4'd9;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd13,6'd26,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd43: Enemy_img = 4'd3;
//6'd34: Enemy_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd30,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd12,6'd27,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd43: Enemy_img = 4'd3;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd13,6'd15,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd11,6'd12,6'd14,6'd16,6'd29,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd44: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd21,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd13,6'd15,6'd18,6'd20,6'd22,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd44: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd24,6'd25,6'd27,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd27,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd37: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd37: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd43,6'd45: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd37: Enemy_img = 4'd13;
//6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//6'd30,6'd31,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd38: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd36,6'd37,6'd39,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd36,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//6'd30,6'd34,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd13;
//6'd31,6'd36,6'd37,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//6'd30,6'd34,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd41: Enemy_img = 4'd13;
//6'd37,6'd38: Enemy_img = 4'd14;
//6'd30,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd13;
//6'd38: Enemy_img = 4'd14;
//6'd31,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd13;
//6'd39: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd13;
//6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd13;
//6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd13;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd28,6'd30,6'd31,6'd32,6'd33,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd3;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd25,6'd28,6'd29,6'd30,6'd31,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd4;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd26,6'd28,6'd30,6'd31,6'd32,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd4;
//6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd33,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd4;
//6'd24,6'd36,6'd37: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd35: Enemy_img = 4'd4;
//6'd24,6'd25,6'd37,6'd38: Enemy_img = 4'd13;
//6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd36,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd4;
//6'd29: Enemy_img = 4'd9;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd24,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd20,6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20: Enemy_img = 4'd3;
//6'd36,6'd37: Enemy_img = 4'd4;
//6'd29: Enemy_img = 4'd9;
//6'd27: Enemy_img = 4'd10;
//6'd21,6'd23,6'd24,6'd25,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21: Enemy_img = 4'd3;
//6'd37,6'd38,6'd39: Enemy_img = 4'd4;
//6'd26: Enemy_img = 4'd9;
//6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd4;
//6'd32: Enemy_img = 4'd9;
//6'd28: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd19,6'd20,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd10;
//6'd20,6'd22,6'd23,6'd24,6'd27,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd42: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd13;
//6'd20,6'd21,6'd27,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd19,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd43: Enemy_img = 4'd3;
//6'd33,6'd35: Enemy_img = 4'd9;
//6'd19,6'd20,6'd21,6'd23,6'd27,6'd30,6'd31,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd18,6'd24,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd44: Enemy_img = 4'd3;
//6'd32: Enemy_img = 4'd9;
//6'd33: Enemy_img = 4'd10;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd30,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd27,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd31,6'd32: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd30,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd17,6'd18: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd16,6'd17,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd27,6'd30,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd26,6'd28,6'd29,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd3;
//6'd37: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46: Enemy_img = 4'd14;
//6'd16,6'd27,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd3;
//6'd38: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd15,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd39: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd15,6'd31,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd44: Enemy_img = 4'd14;
//6'd14,6'd30,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd45: Enemy_img = 4'd14;
//6'd14,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd42,6'd44,6'd45: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd43: Enemy_img = 4'd14;
//6'd13,6'd14,6'd18,6'd19,6'd27,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd3;
//6'd43: Enemy_img = 4'd13;
//6'd14,6'd32,6'd35,6'd36,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd15,6'd16,6'd17,6'd31,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd3;
//6'd44: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd13,6'd15,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd3;
//6'd45: Enemy_img = 4'd13;
//6'd35,6'd41,6'd43,6'd44: Enemy_img = 4'd14;
//6'd33,6'd34,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd13;
//6'd41,6'd44,6'd45: Enemy_img = 4'd14;
//6'd34,6'd35,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd4;
//6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27: Enemy_img = 4'd4;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd4;
//6'd33: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd32,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd4;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd4;
//6'd21: Enemy_img = 4'd13;
//6'd20,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd4;
//6'd24,6'd25: Enemy_img = 4'd9;
//6'd22: Enemy_img = 4'd13;
//6'd20,6'd21,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd38: Enemy_img = 4'd4;
//6'd23: Enemy_img = 4'd9;
//6'd24: Enemy_img = 4'd10;
//6'd20,6'd21,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17,6'd39,6'd40: Enemy_img = 4'd3;
//6'd23,6'd27,6'd28,6'd29: Enemy_img = 4'd9;
//6'd25: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd27: Enemy_img = 4'd10;
//6'd18,6'd19,6'd20,6'd21,6'd25,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd17: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd18: Enemy_img = 4'd3;
//6'd26,6'd31,6'd32: Enemy_img = 4'd9;
//6'd29: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd24,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd17,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd20: Enemy_img = 4'd3;
//6'd26,6'd31: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd18,6'd24,6'd28,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd17,6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd13;
//6'd18,6'd19,6'd28,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd17,6'd21,6'd22,6'd23,6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd9;
//6'd33: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd22,6'd23,6'd24,6'd28,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd16: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22: Enemy_img = 4'd3;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd16: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd25,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd16,6'd24,6'd26,6'd27,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24: Enemy_img = 4'd3;
//6'd37,6'd38: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//6'd15,6'd16,6'd25,6'd26,6'd28,6'd29,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd3;
//6'd39: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd44: Enemy_img = 4'd14;
//6'd15,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd40,6'd41,6'd44: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42: Enemy_img = 4'd14;
//6'd15,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd15,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd3;
//6'd43,6'd44: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd25,6'd26,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd3;
//6'd44,6'd45: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd31,6'd34,6'd35,6'd43: Enemy_img = 4'd14;
//6'd14,6'd23,6'd24,6'd25,6'd26,6'd30,6'd32,6'd33,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd3;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd32,6'd33,6'd34,6'd35,6'd41,6'd44,6'd45: Enemy_img = 4'd14;
//6'd14,6'd20,6'd21,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd3;
//6'd15,6'd16,6'd17,6'd35: Enemy_img = 4'd14;
//6'd14,6'd18,6'd19,6'd33,6'd34,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd15,6'd16: Enemy_img = 4'd14;
//6'd14,6'd17,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd14,6'd15,6'd16: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd14: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42: Enemy_img = 4'd13;
//6'd32,6'd33,6'd43: Enemy_img = 4'd14;
//6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd41: Enemy_img = 4'd13;
//6'd31,6'd32,6'd37,6'd42,6'd43: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd38,6'd40: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd36,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd3;
//6'd39: Enemy_img = 4'd13;
//6'd10,6'd12,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd3;
//6'd38: Enemy_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd4;
//6'd37: Enemy_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd4;
//6'd13,6'd36: Enemy_img = 4'd13;
//6'd11,6'd12,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd4;
//6'd14,6'd15,6'd16,6'd35: Enemy_img = 4'd13;
//6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd4;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd21,6'd34: Enemy_img = 4'd13;
//6'd12,6'd13,6'd20,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24: Enemy_img = 4'd4;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd33: Enemy_img = 4'd13;
//6'd12,6'd13,6'd22,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23: Enemy_img = 4'd4;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd32: Enemy_img = 4'd13;
//6'd13,6'd14,6'd21,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd9;
//6'd16,6'd17,6'd18,6'd19,6'd31: Enemy_img = 4'd13;
//6'd14,6'd15,6'd20,6'd23,6'd24,6'd25,6'd26,6'd27,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd30,6'd31: Enemy_img = 4'd13;
//6'd13,6'd14,6'd15,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd9;
//6'd29: Enemy_img = 4'd10;
//6'd17,6'd18: Enemy_img = 4'd13;
//6'd14,6'd15,6'd16,6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd39,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd20: Enemy_img = 4'd4;
//6'd25,6'd29,6'd30: Enemy_img = 4'd9;
//6'd17: Enemy_img = 4'd13;
//6'd15,6'd16,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd19: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd9;
//6'd27: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28,6'd33,6'd36,6'd37: Enemy_img = 4'd14;
//6'd32,6'd34,6'd35,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd19: Enemy_img = 4'd4;
//6'd26: Enemy_img = 4'd10;
//6'd16,6'd17,6'd18,6'd20,6'd21,6'd24,6'd28,6'd29,6'd30,6'd32: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd18: Enemy_img = 4'd4;
//6'd22,6'd23,6'd27: Enemy_img = 4'd9;
//6'd17,6'd19,6'd20,6'd21,6'd24,6'd31,6'd34,6'd35: Enemy_img = 4'd14;
//6'd32,6'd33,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd25,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd29,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17,6'd18,6'd34,6'd35,6'd36: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd10;
//6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd29,6'd33,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd17,6'd33,6'd34: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd9;
//6'd22: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd29,6'd30,6'd31,6'd35,6'd36: Enemy_img = 4'd14;
//6'd26,6'd28,6'd32,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd3;
//6'd21: Enemy_img = 4'd13;
//6'd17,6'd19,6'd22,6'd23,6'd29,6'd30,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd26,6'd28,6'd31,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd32: Enemy_img = 4'd3;
//6'd20: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd31,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd27,6'd28,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd21,6'd23,6'd24,6'd25,6'd26,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd27,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd3;
//6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd26: Enemy_img = 4'd3;
//6'd23,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24: Enemy_img = 4'd3;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd22,6'd25,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd25,6'd27,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd28,6'd30,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd30,6'd31,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd31,6'd33,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd34,6'd35,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd13;
//6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd13;
//6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd13;
//6'd33,6'd37: Enemy_img = 4'd14;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd28,6'd32,6'd36,6'd37: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd27,6'd32,6'd34,6'd36,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd27,6'd28,6'd33,6'd34,6'd36,6'd37: Enemy_img = 4'd14;
//6'd31,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd33,6'd35,6'd36: Enemy_img = 4'd14;
//6'd31,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd34: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd33,6'd35,6'd36: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd3;
//6'd33: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd3;
//6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd40: Enemy_img = 4'd14;
//6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd4;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd23,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd4;
//6'd32: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd22,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd4;
//6'd32: Enemy_img = 4'd13;
//6'd21,6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39: Enemy_img = 4'd14;
//6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd31: Enemy_img = 4'd13;
//6'd10,6'd12,6'd15,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd9;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd22,6'd23: Enemy_img = 4'd4;
//6'd15,6'd17,6'd18,6'd19,6'd20: Enemy_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd16,6'd21,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd34,6'd37,6'd38: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd29: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Enemy_img = 4'd13;
//6'd10,6'd11,6'd12,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd34: Enemy_img = 4'd14;
//6'd33,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd31: Enemy_img = 4'd9;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Enemy_img = 4'd13;
//6'd11,6'd12,6'd13,6'd21,6'd23,6'd24,6'd25,6'd26,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd27: Enemy_img = 4'd9;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd29: Enemy_img = 4'd13;
//6'd12,6'd13,6'd14,6'd20,6'd21,6'd23,6'd24,6'd25,6'd28,6'd30,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd34,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd27: Enemy_img = 4'd9;
//6'd16,6'd17,6'd18,6'd19,6'd20: Enemy_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd21,6'd23,6'd24,6'd25,6'd31,6'd33,6'd36: Enemy_img = 4'd14;
//6'd34,6'd35,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd21,6'd22: Enemy_img = 4'd4;
//6'd29: Enemy_img = 4'd9;
//6'd28: Enemy_img = 4'd10;
//6'd17,6'd18,6'd19: Enemy_img = 4'd13;
//6'd15,6'd16,6'd20,6'd23,6'd24,6'd25,6'd26,6'd33,6'd34,6'd35,6'd38,6'd39: Enemy_img = 4'd14;
//6'd31,6'd36,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd21: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd9;
//6'd19: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd20,6'd22,6'd23,6'd26,6'd33,6'd34,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd32,6'd35,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd9;
//6'd19,6'd27: Enemy_img = 4'd13;
//6'd17,6'd18,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd33,6'd34,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd31,6'd32,6'd35,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd3;
//6'd21: Enemy_img = 4'd4;
//6'd26: Enemy_img = 4'd9;
//6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd24,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd31,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd3;
//6'd21: Enemy_img = 4'd4;
//6'd27,6'd28,6'd29: Enemy_img = 4'd9;
//6'd19,6'd20,6'd22,6'd23,6'd24,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd30,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd3;
//6'd21: Enemy_img = 4'd4;
//6'd26: Enemy_img = 4'd13;
//6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd30,6'd32,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd31,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd33: Enemy_img = 4'd3;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd32,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd32: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd13;
//6'd22,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd3;
//6'd21,6'd26,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd28,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd3;
//6'd29,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd3;
//6'd41: Enemy_img = 4'd14;
//6'd28,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd30: Enemy_img = 4'd13;
//6'd27,6'd31,6'd33: Enemy_img = 4'd14;
//6'd26,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd27,6'd29,6'd31,6'd32: Enemy_img = 4'd14;
//6'd26,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd27,6'd29,6'd31,6'd32: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd29,6'd31,6'd32: Enemy_img = 4'd14;
//6'd27,6'd34,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd29,6'd31,6'd32,6'd37: Enemy_img = 4'd14;
//6'd27,6'd34,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd29,6'd31,6'd32,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd39: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd39: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd39: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd39: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd21,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd21,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd13;
//6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd31,6'd32,6'd34,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd35,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd9;
//6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd33,6'd35,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd29,6'd31,6'd32: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd27,6'd34,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd35,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd33,6'd34,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd21,6'd30: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd22,6'd24,6'd25,6'd26,6'd27,6'd29,6'd31,6'd32,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd37,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd9;
//6'd19,6'd20,6'd21: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd22,6'd24,6'd25,6'd26,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd33,6'd37,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd29,6'd31,6'd32: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd18,6'd19,6'd20,6'd21: Enemy_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd22,6'd24,6'd25,6'd26,6'd27,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd34,6'd37,6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd4;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Enemy_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd33,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd34,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd28,6'd33,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd4;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd30: Enemy_img = 4'd13;
//default: Enemy_img = 4'd14;
//6'd34,6'd35,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd4;
//6'd28: Enemy_img = 4'd9;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Enemy_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd23,6'd25,6'd26,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd33,6'd35,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd4;
//6'd29,6'd31,6'd32: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd19,6'd20,6'd21,6'd22: Enemy_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd23,6'd25,6'd26,6'd27,6'd34,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd35,6'd36,6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd4;
//6'd22: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd26,6'd27,6'd28,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd4;
//6'd30: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd35: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd24,6'd25,6'd27,6'd28,6'd31,6'd34: Enemy_img = 4'd14;
//6'd33,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd35: Enemy_img = 4'd3;
//6'd27: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd13;
//6'd25: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd13;
//6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd13;
//6'd26: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd27: Enemy_img = 4'd14;
//6'd30,6'd31,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd26: Enemy_img = 4'd13;
//6'd27,6'd28: Enemy_img = 4'd14;
//6'd30,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd13;
//6'd23,6'd25,6'd27,6'd28,6'd29,6'd34: Enemy_img = 4'd14;
//6'd22,6'd31,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd13;
//6'd23,6'd24,6'd26,6'd28,6'd29,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd22,6'd31,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd27: Enemy_img = 4'd13;
//6'd24,6'd26,6'd28,6'd29,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd28: Enemy_img = 4'd13;
//6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36: Enemy_img = 4'd14;
//6'd24,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd28: Enemy_img = 4'd13;
//6'd20,6'd22,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd28: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd39: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd35,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd39: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd44: Enemy_img = 4'd14;
//6'd35,6'd43,6'd45,6'd47,6'd50,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd39: Enemy_img = 4'd3;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd33,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd52: Enemy_img = 4'd14;
//6'd34,6'd36,6'd49,6'd51,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd39,6'd40: Enemy_img = 4'd3;
//6'd31: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd35,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd29,6'd32,6'd33: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd22,6'd39,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd31: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd27,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd22,6'd39,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd23: Enemy_img = 4'd4;
//6'd32: Enemy_img = 4'd13;
//6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd35,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd3;
//6'd24,6'd25: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd9;
//6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd31,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd37,6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd4;
//6'd31,6'd34: Enemy_img = 4'd9;
//6'd33: Enemy_img = 4'd10;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd36,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd26: Enemy_img = 4'd4;
//6'd32: Enemy_img = 4'd9;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd36,6'd40,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd39,6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd4;
//6'd24,6'd34: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd37,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd27,6'd28: Enemy_img = 4'd4;
//6'd36: Enemy_img = 4'd9;
//6'd23,6'd24: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd25,6'd26,6'd29,6'd30,6'd31,6'd38,6'd39,6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd28: Enemy_img = 4'd4;
//6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd35: Enemy_img = 4'd10;
//6'd23,6'd24,6'd25: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd26,6'd27,6'd29,6'd30,6'd38,6'd39,6'd40,6'd42: Enemy_img = 4'd14;
//6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd28,6'd29: Enemy_img = 4'd4;
//6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd27,6'd30,6'd31,6'd32,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd4;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd35: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd30: Enemy_img = 4'd4;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd36: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd4;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd36: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd26,6'd27,6'd29,6'd30,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd3;
//6'd31: Enemy_img = 4'd4;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd3;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd31,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd20: Enemy_img = 4'd14;
//6'd25,6'd26,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19: Enemy_img = 4'd13;
//6'd20,6'd21,6'd24: Enemy_img = 4'd14;
//6'd25,6'd26,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd3;
//6'd20: Enemy_img = 4'd13;
//6'd21,6'd22,6'd24,6'd30: Enemy_img = 4'd14;
//6'd26,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd3;
//6'd21: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd27,6'd50,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd3;
//6'd22: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd29,6'd30,6'd33,6'd51: Enemy_img = 4'd14;
//6'd31,6'd32,6'd34,6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd3;
//6'd20,6'd21,6'd23: Enemy_img = 4'd13;
//6'd22,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd34,6'd35,6'd46,6'd47,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd13;
//6'd20,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd19,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd25: Enemy_img = 4'd13;
//6'd21,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd19,6'd20,6'd35,6'd36,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd26: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd22,6'd34,6'd35,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd3;
//6'd27: Enemy_img = 4'd13;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd34,6'd35,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd3;
//6'd28: Enemy_img = 4'd13;
//6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd35,6'd36,6'd38,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd3;
//6'd29: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd35,6'd38,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd34,6'd36,6'd37,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd40,6'd48,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd33,6'd34: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd35,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd42: Enemy_img = 4'd3;
//6'd33: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd35,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd43: Enemy_img = 4'd3;
//6'd30,6'd32: Enemy_img = 4'd9;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35,6'd38,6'd42,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd43: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd38,6'd44,6'd45: Enemy_img = 4'd14;
//6'd41,6'd42,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44: Enemy_img = 4'd3;
//6'd24: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd10;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd38,6'd41,6'd42,6'd43,6'd45: Enemy_img = 4'd14;
//6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd4;
//6'd33: Enemy_img = 4'd9;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd37,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd23,6'd24,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd3;
//6'd26,6'd27,6'd28: Enemy_img = 4'd4;
//6'd39: Enemy_img = 4'd9;
//6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45: Enemy_img = 4'd3;
//6'd28,6'd29: Enemy_img = 4'd4;
//6'd36: Enemy_img = 4'd9;
//6'd38: Enemy_img = 4'd10;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42,6'd44: Enemy_img = 4'd14;
//6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd4;
//6'd36: Enemy_img = 4'd9;
//6'd39: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41: Enemy_img = 4'd14;
//6'd43,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd32: Enemy_img = 4'd4;
//6'd27,6'd28,6'd40: Enemy_img = 4'd13;
//6'd25,6'd26,6'd29,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd4;
//6'd28,6'd29,6'd41: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd4;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd13;
//6'd25,6'd26,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd3;
//6'd36: Enemy_img = 4'd4;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd25,6'd26,6'd33,6'd34,6'd35,6'd37,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd3;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd34,6'd35,6'd36,6'd37,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd13;
//6'd24,6'd25,6'd32,6'd33,6'd34,6'd35,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd13;
//6'd24,6'd25,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd13;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd24: Enemy_img = 4'd14;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd14;
//6'd46,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd14;
//6'd45,6'd46,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd44,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd43,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd26,6'd41,6'd43,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd3;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd27,6'd28,6'd39,6'd40,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd3;
//6'd26,6'd27,6'd28,6'd30,6'd31,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd22,6'd23,6'd29,6'd36,6'd37,6'd38,6'd40,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd3;
//6'd27,6'd28,6'd29,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd37,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd3;
//6'd17,6'd21,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd29,6'd34,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd3;
//6'd17: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd22,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd34,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd3;
//6'd18,6'd19: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd33,6'd34,6'd38,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd3;
//6'd20,6'd21,6'd22: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd36,6'd38,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd37,6'd39,6'd40,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43: Enemy_img = 4'd3;
//6'd23,6'd24: Enemy_img = 4'd13;
//6'd21,6'd22,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd36,6'd37,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44: Enemy_img = 4'd3;
//6'd25,6'd26,6'd27: Enemy_img = 4'd13;
//6'd19,6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd45,6'd46: Enemy_img = 4'd14;
//6'd34,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45: Enemy_img = 4'd3;
//6'd27,6'd28,6'd29: Enemy_img = 4'd13;
//6'd20,6'd21,6'd25,6'd26,6'd30,6'd31,6'd32,6'd33,6'd36,6'd41,6'd43,6'd46,6'd47: Enemy_img = 4'd14;
//6'd19,6'd39,6'd40,6'd42,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd3;
//6'd35: Enemy_img = 4'd9;
//6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd33,6'd37,6'd44,6'd45: Enemy_img = 4'd14;
//6'd19,6'd20,6'd22,6'd23,6'd38,6'd40,6'd41,6'd43,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd3;
//6'd39: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd10;
//6'd32: Enemy_img = 4'd13;
//6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd36,6'd40,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd3;
//6'd34,6'd38,6'd42: Enemy_img = 4'd9;
//6'd36: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd40,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd42: Enemy_img = 4'd9;
//6'd38: Enemy_img = 4'd10;
//6'd20,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd36,6'd40,6'd44,6'd45: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd42: Enemy_img = 4'd9;
//6'd40: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd9;
//6'd43,6'd44: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd3;
//6'd40: Enemy_img = 4'd9;
//6'd44,6'd45: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd3;
//6'd27: Enemy_img = 4'd4;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd4;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd4;
//6'd29,6'd30,6'd31,6'd32,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd3;
//6'd38,6'd39,6'd41,6'd42,6'd43: Enemy_img = 4'd4;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd37: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd31,6'd32,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd13;
//6'd32,6'd33,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd13;
//6'd31,6'd32,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd32,6'd33,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd13;
//6'd32,6'd33,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd14;
//6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd14;
//6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd39,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd39,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd38,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd38,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd37,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd36,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd35,6'd36,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd34,6'd35,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd33,6'd34,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd3;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd3;
//6'd27,6'd28,6'd33,6'd34,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd3;
//6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd28,6'd32,6'd36,6'd37,6'd38,6'd39,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46: Enemy_img = 4'd3;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd27,6'd32,6'd36,6'd43,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd20,6'd21,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd39,6'd40,6'd41,6'd48,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd36,6'd40,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd34,6'd38,6'd42,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd39,6'd43: Enemy_img = 4'd9;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd41,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd39,6'd43: Enemy_img = 4'd9;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd41,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd39,6'd43: Enemy_img = 4'd10;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd41,6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd39,6'd43: Enemy_img = 4'd9;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd41,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd38,6'd42: Enemy_img = 4'd9;
//6'd20: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd36,6'd40,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd20,6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46: Enemy_img = 4'd4;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd4;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd4;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd4;
//6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42: Enemy_img = 4'd13;
//6'd38,6'd39,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd13;
//6'd39,6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_0 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd14;
//6'd32,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd14;
//6'd33,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd32,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd33,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd32,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd32,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd31,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd31,6'd32,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd31,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd3;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41: Enemy_img = 4'd14;
//6'd30,6'd31,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd3;
//6'd32,6'd33,6'd40,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd30,6'd31,6'd41,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd3;
//6'd37,6'd38,6'd39,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd35,6'd36,6'd40,6'd41,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd3;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd29,6'd30,6'd34,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd3;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd38,6'd39,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42: Enemy_img = 4'd9;
//6'd46,6'd47: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd35,6'd36,6'd39,6'd40,6'd44,6'd45: Enemy_img = 4'd14;
//6'd30,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd9;
//6'd43: Enemy_img = 4'd10;
//6'd45: Enemy_img = 4'd13;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd41,6'd46: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd26,6'd31,6'd32,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd43: Enemy_img = 4'd9;
//6'd41: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd37,6'd45,6'd46,6'd47,6'd49,6'd50: Enemy_img = 4'd14;
//6'd21,6'd26,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd3;
//6'd35,6'd43: Enemy_img = 4'd9;
//6'd39: Enemy_img = 4'd10;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd41,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd3;
//6'd35,6'd40,6'd43: Enemy_img = 4'd9;
//6'd37: Enemy_img = 4'd13;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd41,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd4;
//6'd36,6'd39: Enemy_img = 4'd9;
//6'd33,6'd34: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd38,6'd41,6'd42,6'd44,6'd45,6'd46,6'd49: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd4;
//6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd4;
//6'd35: Enemy_img = 4'd9;
//6'd29,6'd30: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd20: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44: Enemy_img = 4'd4;
//6'd26,6'd27,6'd28,6'd47: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42: Enemy_img = 4'd4;
//6'd24,6'd25,6'd45,6'd46: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd4;
//6'd21,6'd22,6'd23,6'd44,6'd45,6'd46: Enemy_img = 4'd13;
//6'd19,6'd20,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd4;
//6'd19,6'd20,6'd21,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//6'd18,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd4;
//6'd18,6'd22,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd48,6'd49: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd4;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//6'd23,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd40,6'd41,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd3;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49: Enemy_img = 4'd14;
//6'd23,6'd24,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd3;
//6'd45,6'd46,6'd47: Enemy_img = 4'd13;
//6'd28,6'd29,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd27,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//2'd1: begin
//case(angle)
//// Enemy_type_1 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd30,6'd31,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd28,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd13;
//6'd26,6'd37,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd2;
//6'd40,6'd41: Enemy_img = 4'd13;
//6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd1;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd2;
//6'd22,6'd26,6'd27,6'd28,6'd29,6'd30,6'd40,6'd41: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd37: Enemy_img = 4'd2;
//6'd21,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd2;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd26,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd10;
//6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd9;
//6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd26,6'd27,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd21,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd37: Enemy_img = 4'd1;
//6'd21: Enemy_img = 4'd14;
//6'd22,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd1;
//6'd22,6'd40,6'd41: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd1;
//6'd40,6'd41: Enemy_img = 4'd13;
//6'd23: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd1;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41: Enemy_img = 4'd14;
//6'd26,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd28,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd30,6'd31,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd28,6'd29,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd33: Enemy_img = 4'd13;
//6'd27,6'd30,6'd31,6'd32,6'd34: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd33,6'd34,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd2;
//6'd28,6'd29,6'd36,6'd37: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd2;
//6'd26,6'd27,6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd25,6'd28,6'd29,6'd33,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd2;
//6'd28,6'd29,6'd30: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd2;
//6'd26,6'd27: Enemy_img = 4'd13;
//6'd24,6'd25,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd2;
//6'd24,6'd25: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd2;
//6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd2;
//6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd21,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd2;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd21,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd36,6'd37: Enemy_img = 4'd14;
//6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd20,6'd25,6'd26,6'd27,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd9;
//6'd29: Enemy_img = 4'd10;
//6'd31: Enemy_img = 4'd13;
//6'd20,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd28: Enemy_img = 4'd10;
//6'd26: Enemy_img = 4'd13;
//6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd1;
//6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd25,6'd26,6'd42: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd1;
//6'd41: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd32,6'd33,6'd34,6'd42: Enemy_img = 4'd14;
//6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd39: Enemy_img = 4'd1;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd1;
//6'd29,6'd37,6'd38: Enemy_img = 4'd14;
//6'd28,6'd35,6'd36,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd1;
//6'd35,6'd36,6'd40: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd38,6'd39: Enemy_img = 4'd14;
//6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd33,6'd34,6'd38,6'd39,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd33,6'd34,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd36,6'd37: Enemy_img = 4'd14;
//6'd31,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd25,6'd26,6'd28: Enemy_img = 4'd14;
//6'd19,6'd20,6'd21,6'd23,6'd24,6'd27,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd1;
//6'd21,6'd22,6'd24,6'd25,6'd27: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd23,6'd26,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd1;
//6'd20,6'd21,6'd23,6'd24,6'd26: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19,6'd22,6'd25,6'd27,6'd28,6'd29,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd1;
//6'd19,6'd20,6'd22,6'd23,6'd25,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd16,6'd17,6'd18,6'd21,6'd24,6'd26,6'd27,6'd28,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd22,6'd24,6'd30,6'd31,6'd32,6'd34,6'd35: Enemy_img = 4'd14;
//6'd15,6'd16,6'd17,6'd20,6'd23,6'd25,6'd26,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd32,6'd33: Enemy_img = 4'd9;
//6'd35: Enemy_img = 4'd13;
//6'd18,6'd20,6'd21,6'd23,6'd29,6'd36: Enemy_img = 4'd14;
//6'd14,6'd15,6'd16,6'd17,6'd19,6'd22,6'd24,6'd25,6'd27,6'd28,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd31,6'd32,6'd33: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd10;
//6'd20,6'd28,6'd29,6'd36: Enemy_img = 4'd14;
//6'd14,6'd16,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd24: Enemy_img = 4'd1;
//6'd38: Enemy_img = 4'd2;
//6'd31,6'd32: Enemy_img = 4'd9;
//6'd33: Enemy_img = 4'd10;
//6'd27,6'd28,6'd29,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd25,6'd26,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24: Enemy_img = 4'd1;
//6'd37,6'd38: Enemy_img = 4'd2;
//6'd33: Enemy_img = 4'd9;
//6'd20,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36,6'd39: Enemy_img = 4'd14;
//6'd25,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd1;
//6'd36,6'd37: Enemy_img = 4'd2;
//6'd20,6'd31: Enemy_img = 4'd13;
//6'd19,6'd28,6'd29,6'd30,6'd35,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd2;
//6'd20,6'd30: Enemy_img = 4'd13;
//6'd21,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd2;
//6'd29,6'd39: Enemy_img = 4'd13;
//6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd2;
//6'd28,6'd38: Enemy_img = 4'd13;
//6'd26,6'd27,6'd29,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd2;
//6'd27,6'd37,6'd39: Enemy_img = 4'd13;
//6'd26,6'd28,6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd33: Enemy_img = 4'd2;
//6'd36,6'd38,6'd39: Enemy_img = 4'd13;
//6'd31,6'd32,6'd34,6'd35,6'd37,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd2;
//6'd35,6'd37,6'd38: Enemy_img = 4'd13;
//6'd33,6'd34,6'd36,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd2;
//6'd34,6'd36,6'd37: Enemy_img = 4'd13;
//6'd32,6'd33,6'd35,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd2;
//6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd2;
//6'd34,6'd35,6'd37,6'd38: Enemy_img = 4'd13;
//6'd29,6'd33,6'd36,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd33,6'd34,6'd36,6'd37: Enemy_img = 4'd13;
//6'd32,6'd35,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd13;
//6'd30,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd13;
//6'd32,6'd33,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd14;
//6'd27,6'd28,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd1;
//6'd26,6'd39: Enemy_img = 4'd14;
//6'd24,6'd25,6'd27,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd1;
//6'd26,6'd32,6'd33,6'd40: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd30,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd1;
//6'd34: Enemy_img = 4'd13;
//6'd23,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd40: Enemy_img = 4'd14;
//6'd21,6'd22,6'd24,6'd26,6'd27,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd1;
//6'd23,6'd25,6'd29,6'd30,6'd34: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd24,6'd26,6'd27,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd2;
//6'd31,6'd32: Enemy_img = 4'd9;
//6'd20,6'd22,6'd24,6'd28,6'd29,6'd34,6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd30,6'd31,6'd33: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd20,6'd22,6'd24,6'd28,6'd35,6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd30,6'd31,6'd33: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd39: Enemy_img = 4'd13;
//6'd19,6'd21,6'd23,6'd24,6'd28,6'd35,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd17,6'd18,6'd20,6'd22,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd33: Enemy_img = 4'd9;
//6'd39: Enemy_img = 4'd13;
//6'd19,6'd21,6'd23,6'd27,6'd28,6'd29,6'd31,6'd35,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//6'd17,6'd18,6'd20,6'd22,6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd31,6'd38,6'd39,6'd41: Enemy_img = 4'd13;
//6'd18,6'd21,6'd23,6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd37,6'd40: Enemy_img = 4'd14;
//6'd16,6'd17,6'd19,6'd20,6'd22,6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd31,6'd38,6'd40: Enemy_img = 4'd13;
//6'd18,6'd20,6'd26,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//6'd16,6'd17,6'd19,6'd21,6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd30,6'd38,6'd40: Enemy_img = 4'd13;
//6'd18,6'd20,6'd26,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//6'd16,6'd17,6'd19,6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd1;
//6'd35: Enemy_img = 4'd2;
//6'd30,6'd37,6'd39: Enemy_img = 4'd13;
//6'd20,6'd21,6'd28,6'd29,6'd31,6'd33,6'd34,6'd36,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd2;
//6'd22,6'd29,6'd30,6'd37,6'd39,6'd41: Enemy_img = 4'd13;
//6'd21,6'd28,6'd31,6'd33,6'd34,6'd36,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//6'd17: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd2;
//6'd22,6'd29,6'd36,6'd39,6'd41: Enemy_img = 4'd13;
//6'd21,6'd23,6'd28,6'd35,6'd37,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd2;
//6'd36,6'd38,6'd40: Enemy_img = 4'd13;
//6'd28,6'd35,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd2;
//6'd38,6'd40: Enemy_img = 4'd13;
//6'd36,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd39,6'd40: Enemy_img = 4'd13;
//6'd36,6'd38,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd39: Enemy_img = 4'd13;
//6'd33,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd39: Enemy_img = 4'd13;
//6'd34,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd36: Enemy_img = 4'd14;
//6'd28,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd37: Enemy_img = 4'd14;
//6'd27,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd14;
//6'd26,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd13;
//6'd31: Enemy_img = 4'd14;
//6'd25,6'd26,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd32: Enemy_img = 4'd13;
//6'd30,6'd31,6'd33,6'd35,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd39: Enemy_img = 4'd13;
//6'd24,6'd29,6'd30,6'd33,6'd34,6'd35,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd23,6'd25,6'd26,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd31: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd39: Enemy_img = 4'd13;
//6'd24,6'd28,6'd29,6'd34,6'd35,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//6'd22,6'd23,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd30,6'd31,6'd33: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd39,6'd41: Enemy_img = 4'd13;
//6'd22,6'd24,6'd28,6'd35,6'd37,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//6'd21,6'd23,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd30,6'd31,6'd33: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd39,6'd41: Enemy_img = 4'd13;
//6'd22,6'd24,6'd28,6'd35,6'd37,6'd38,6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd30,6'd33: Enemy_img = 4'd9;
//6'd39,6'd41: Enemy_img = 4'd13;
//6'd22,6'd24,6'd28,6'd35,6'd36,6'd38,6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd32,6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd28,6'd29,6'd31,6'd34,6'd35,6'd36,6'd38,6'd40,6'd42,6'd44: Enemy_img = 4'd14;
//6'd19,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd32,6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd38,6'd40,6'd42,6'd44: Enemy_img = 4'd14;
//6'd19,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd32,6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd32,6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd28,6'd30,6'd31,6'd33,6'd35,6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd32,6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd28,6'd30,6'd31,6'd33,6'd35,6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28: Enemy_img = 4'd1;
//6'd35,6'd36,6'd37: Enemy_img = 4'd2;
//6'd32,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd31,6'd33,6'd38,6'd39,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd23,6'd24,6'd25,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd37: Enemy_img = 4'd1;
//6'd38,6'd39: Enemy_img = 4'd2;
//6'd32,6'd41,6'd43: Enemy_img = 4'd13;
//6'd20,6'd22,6'd31,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd43: Enemy_img = 4'd13;
//6'd20,6'd23,6'd31,6'd41,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd21,6'd22,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd13;
//6'd24,6'd26,6'd37,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd13;
//6'd24,6'd26,6'd37,6'd39,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd45: Enemy_img = 4'd14;
//6'd18,6'd20: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd14;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd14;
//6'd24,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd2;
//6'd36: Enemy_img = 4'd13;
//6'd23,6'd34,6'd35,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd2;
//6'd29,6'd36: Enemy_img = 4'd13;
//6'd22,6'd32,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd2;
//6'd29,6'd30,6'd37,6'd39: Enemy_img = 4'd13;
//6'd22,6'd28,6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd2;
//6'd37,6'd39: Enemy_img = 4'd13;
//6'd27,6'd28,6'd32,6'd33,6'd35,6'd36,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd35: Enemy_img = 4'd2;
//6'd31: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd38,6'd40,6'd42: Enemy_img = 4'd13;
//6'd27,6'd28,6'd33,6'd34,6'd36,6'd37,6'd39,6'd41,6'd43,6'd44: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd29,6'd30,6'd32: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd10;
//6'd38,6'd40,6'd42: Enemy_img = 4'd13;
//6'd26,6'd27,6'd34,6'd35,6'd37,6'd39,6'd41,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd2;
//6'd29,6'd30,6'd32: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd10;
//6'd38,6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd23,6'd27,6'd34,6'd35,6'd37,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd22,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd39,6'd41,6'd43: Enemy_img = 4'd13;
//6'd23,6'd27,6'd31,6'd33,6'd34,6'd35,6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd14;
//6'd21,6'd22,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37: Enemy_img = 4'd2;
//6'd32,6'd39,6'd41,6'd44: Enemy_img = 4'd13;
//6'd21,6'd23,6'd24,6'd28,6'd31,6'd33,6'd34,6'd35,6'd36,6'd38,6'd40,6'd42,6'd43,6'd45,6'd46: Enemy_img = 4'd14;
//6'd22,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37,6'd38: Enemy_img = 4'd2;
//6'd32,6'd42,6'd44: Enemy_img = 4'd13;
//6'd22,6'd24,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd36,6'd39,6'd40,6'd41,6'd43,6'd45,6'd46: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd2;
//6'd33,6'd44: Enemy_img = 4'd13;
//6'd22,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd36,6'd41,6'd42,6'd43,6'd45,6'd46: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd39: Enemy_img = 4'd2;
//6'd33: Enemy_img = 4'd13;
//6'd23,6'd25,6'd29,6'd31,6'd32,6'd34,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd24,6'd26,6'd28,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd34,6'd40: Enemy_img = 4'd13;
//6'd21,6'd23,6'd25,6'd29,6'd32,6'd33,6'd41,6'd45: Enemy_img = 4'd14;
//6'd20,6'd22,6'd24,6'd26,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd1;
//6'd34,6'd40: Enemy_img = 4'd13;
//6'd21,6'd23,6'd26,6'd33,6'd39,6'd41: Enemy_img = 4'd14;
//6'd20,6'd22,6'd24,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd1;
//6'd34: Enemy_img = 4'd13;
//6'd22,6'd24,6'd26: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd25,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd1;
//6'd22,6'd24: Enemy_img = 4'd14;
//6'd20,6'd21,6'd23,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd25: Enemy_img = 4'd14;
//6'd20,6'd21,6'd24,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd13;
//6'd23,6'd29: Enemy_img = 4'd14;
//6'd21,6'd22,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd13;
//6'd23,6'd28: Enemy_img = 4'd14;
//6'd21,6'd22,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd36,6'd37,6'd40: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd35,6'd38,6'd39,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd2;
//6'd35,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd36,6'd39,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd2;
//6'd36,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd13;
//6'd30,6'd33,6'd34,6'd35,6'd37,6'd40,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd2;
//6'd27,6'd37,6'd39,6'd40,6'd42,6'd43: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd38,6'd41,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd2;
//6'd28,6'd38,6'd40,6'd41,6'd43,6'd44: Enemy_img = 4'd13;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd36,6'd37,6'd39,6'd42,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd2;
//6'd29: Enemy_img = 4'd10;
//6'd39,6'd41,6'd42,6'd44: Enemy_img = 4'd13;
//6'd26,6'd27,6'd33,6'd34,6'd35,6'd37,6'd38,6'd40,6'd43,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd2;
//6'd28,6'd29,6'd31: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd42: Enemy_img = 4'd13;
//6'd26,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd48: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd1;
//6'd38,6'd41: Enemy_img = 4'd2;
//6'd28,6'd29,6'd30,6'd32: Enemy_img = 4'd9;
//6'd26,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd21,6'd22,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd1;
//6'd38,6'd39,6'd40: Enemy_img = 4'd2;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd13;
//6'd26,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd1;
//6'd37,6'd38: Enemy_img = 4'd2;
//6'd30: Enemy_img = 4'd9;
//6'd33,6'd42: Enemy_img = 4'd13;
//6'd27,6'd31,6'd32,6'd34,6'd43: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd1;
//6'd34,6'd42: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd41: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd35: Enemy_img = 4'd13;
//6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36: Enemy_img = 4'd14;
//6'd22,6'd24,6'd25,6'd26,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd1;
//6'd36: Enemy_img = 4'd13;
//6'd24,6'd30,6'd31,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd22,6'd23,6'd25,6'd26,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd1;
//6'd23,6'd25,6'd31,6'd35,6'd36: Enemy_img = 4'd14;
//6'd22,6'd24,6'd26,6'd27,6'd29,6'd30,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd32: Enemy_img = 4'd1;
//6'd23,6'd24,6'd26: Enemy_img = 4'd14;
//6'd22,6'd25,6'd27,6'd28,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd1;
//6'd24,6'd25,6'd27: Enemy_img = 4'd14;
//6'd22,6'd23,6'd26,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd1;
//6'd25,6'd26,6'd28: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd27,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd1;
//6'd23,6'd24,6'd26,6'd27: Enemy_img = 4'd14;
//6'd25,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd1;
//6'd24,6'd25,6'd27,6'd28,6'd33: Enemy_img = 4'd14;
//6'd23,6'd26,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd25,6'd26,6'd28,6'd29,6'd31: Enemy_img = 4'd14;
//6'd23,6'd24,6'd27,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd32: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd36,6'd37: Enemy_img = 4'd13;
//6'd31,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd38,6'd39,6'd40: Enemy_img = 4'd13;
//6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42: Enemy_img = 4'd13;
//6'd23,6'd24,6'd28,6'd29,6'd33,6'd34,6'd38,6'd39,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd38,6'd39: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd23,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd2;
//6'd35,6'd36,6'd40: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd2;
//6'd37,6'd38: Enemy_img = 4'd13;
//6'd28,6'd29,6'd35,6'd36,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd39: Enemy_img = 4'd2;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd2;
//6'd26,6'd41: Enemy_img = 4'd13;
//6'd27,6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd2;
//6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd42: Enemy_img = 4'd13;
//6'd25,6'd26,6'd33,6'd34,6'd35,6'd36,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd2;
//6'd28: Enemy_img = 4'd9;
//6'd29,6'd30: Enemy_img = 4'd10;
//6'd25,6'd26,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd9;
//6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd20,6'd26,6'd34,6'd35: Enemy_img = 4'd14;
//6'd21: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd34,6'd35,6'd36: Enemy_img = 4'd13;
//6'd20,6'd26,6'd27,6'd32,6'd33: Enemy_img = 4'd14;
//6'd21,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd1;
//6'd36,6'd37: Enemy_img = 4'd13;
//6'd21,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd1;
//6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd1;
//6'd24,6'd25,6'd33,6'd34: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd1;
//6'd26,6'd27: Enemy_img = 4'd14;
//6'd24,6'd25,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd1;
//6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd1;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd37: Enemy_img = 4'd14;
//6'd25,6'd28,6'd29,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd1;
//6'd36,6'd37: Enemy_img = 4'd13;
//6'd28,6'd29: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd27,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd14;
//6'd28,6'd29,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd28,6'd29,6'd32,6'd33: Enemy_img = 4'd13;
//6'd23,6'd24,6'd27,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd2;
//6'd24,6'd25,6'd27,6'd28: Enemy_img = 4'd13;
//6'd23,6'd26,6'd29,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd2;
//6'd23,6'd24,6'd26,6'd27: Enemy_img = 4'd13;
//6'd25,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd2;
//6'd25,6'd26,6'd28: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd27,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd2;
//6'd24,6'd25,6'd27: Enemy_img = 4'd13;
//6'd22,6'd23,6'd26,6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd32: Enemy_img = 4'd2;
//6'd23,6'd24,6'd26: Enemy_img = 4'd13;
//6'd22,6'd25,6'd27,6'd28,6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd2;
//6'd23,6'd25,6'd35,6'd36: Enemy_img = 4'd13;
//6'd22,6'd24,6'd26,6'd27,6'd29,6'd30,6'd31,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd2;
//6'd24,6'd34,6'd35: Enemy_img = 4'd13;
//6'd22,6'd23,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd33,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd2;
//6'd23,6'd33,6'd34: Enemy_img = 4'd13;
//6'd22,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd2;
//6'd32,6'd33,6'd42: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd1;
//6'd25,6'd26: Enemy_img = 4'd2;
//6'd30: Enemy_img = 4'd9;
//6'd31,6'd32,6'd42: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd27,6'd33,6'd34,6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40: Enemy_img = 4'd1;
//6'd24,6'd25: Enemy_img = 4'd2;
//6'd29: Enemy_img = 4'd9;
//6'd23,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd21,6'd22,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd41: Enemy_img = 4'd1;
//6'd24: Enemy_img = 4'd2;
//6'd31,6'd32: Enemy_img = 4'd9;
//6'd29,6'd30: Enemy_img = 4'd10;
//6'd25,6'd26,6'd27,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd21,6'd22,6'd36,6'd37,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd30,6'd31: Enemy_img = 4'd9;
//6'd28,6'd29: Enemy_img = 4'd10;
//6'd26,6'd33,6'd34,6'd42: Enemy_img = 4'd14;
//6'd21,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd27: Enemy_img = 4'd13;
//6'd26,6'd33,6'd39,6'd41,6'd42,6'd44: Enemy_img = 4'd14;
//6'd21,6'd34,6'd35,6'd37,6'd38,6'd40,6'd43,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd1;
//6'd26,6'd27: Enemy_img = 4'd13;
//6'd28,6'd30,6'd31,6'd32,6'd38,6'd40,6'd41,6'd43,6'd44: Enemy_img = 4'd14;
//6'd21,6'd36,6'd37,6'd39,6'd42,6'd45,6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd1;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd39,6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//6'd21,6'd34,6'd35,6'd36,6'd38,6'd41,6'd44,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd1;
//6'd36,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//6'd30,6'd33,6'd34,6'd35,6'd37,6'd40,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd1;
//6'd35,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd36,6'd39,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd36,6'd37,6'd40: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd35,6'd38,6'd39,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd29: Enemy_img = 4'd13;
//6'd21,6'd22,6'd24,6'd25,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd28: Enemy_img = 4'd13;
//6'd21,6'd22,6'd24,6'd25,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd25: Enemy_img = 4'd13;
//6'd20,6'd21,6'd24,6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd2;
//6'd22,6'd24: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd2;
//6'd22,6'd24,6'd26: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd27,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd2;
//6'd21,6'd23,6'd26,6'd33,6'd40: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd25,6'd27,6'd34,6'd39,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd2;
//6'd21,6'd23,6'd25,6'd32,6'd33,6'd40: Enemy_img = 4'd13;
//6'd20,6'd22,6'd24,6'd26,6'd28,6'd29,6'd34,6'd41: Enemy_img = 4'd14;
//6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd23,6'd25,6'd32: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd24,6'd26,6'd28,6'd29,6'd31,6'd33,6'd34,6'd41,6'd42: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd22,6'd24,6'd32: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd36,6'd42,6'd44: Enemy_img = 4'd14;
//6'd41,6'd43,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd22,6'd24,6'd31: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd36,6'd42,6'd44: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd43,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd21,6'd23,6'd24,6'd31: Enemy_img = 4'd13;
//6'd22,6'd25,6'd27,6'd28,6'd32,6'd33,6'd34,6'd35,6'd39,6'd41,6'd44: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd43,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd29: Enemy_img = 4'd9;
//6'd23: Enemy_img = 4'd13;
//6'd21,6'd22,6'd24,6'd25,6'd27,6'd34,6'd35,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd29,6'd31,6'd32: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd23: Enemy_img = 4'd13;
//6'd22,6'd24,6'd25,6'd27,6'd34,6'd38,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd35,6'd37,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd25: Enemy_img = 4'd2;
//6'd29,6'd31,6'd32: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd34,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//6'd35,6'd37,6'd39,6'd41,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd2;
//6'd30,6'd31: Enemy_img = 4'd9;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd33,6'd34,6'd38,6'd40,6'd42: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd39,6'd41,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd1;
//6'd28,6'd32,6'd33,6'd37,6'd39: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd35,6'd36,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd1;
//6'd28: Enemy_img = 4'd13;
//6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd39: Enemy_img = 4'd14;
//6'd23,6'd35,6'd36,6'd38,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd1;
//6'd22,6'd29,6'd30,6'd36: Enemy_img = 4'd14;
//6'd23,6'd32,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd1;
//6'd23,6'd36: Enemy_img = 4'd14;
//6'd34,6'd35,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd14;
//6'd24,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd14;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd18,6'd20: Enemy_img = 4'd14;
//6'd43,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd24,6'd26,6'd37,6'd39: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd24,6'd26,6'd37,6'd39: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd22,6'd32,6'd40,6'd43: Enemy_img = 4'd14;
//6'd23,6'd41,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd37,6'd38,6'd39: Enemy_img = 4'd1;
//6'd24,6'd25: Enemy_img = 4'd2;
//6'd20,6'd22,6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd23,6'd32,6'd41,6'd43: Enemy_img = 4'd14;
//6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd1;
//6'd26,6'd27,6'd28: Enemy_img = 4'd2;
//6'd20,6'd22,6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd23,6'd24,6'd25,6'd30,6'd32,6'd41,6'd43: Enemy_img = 4'd14;
//6'd33,6'd38,6'd39,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd20,6'd22,6'd24,6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd27,6'd28,6'd30,6'd32,6'd33,6'd35,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd20,6'd22,6'd24,6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd27,6'd28,6'd30,6'd32,6'd33,6'd35,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd20,6'd22,6'd24,6'd31: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd20,6'd22,6'd24,6'd31: Enemy_img = 4'd13;
//6'd19,6'd21,6'd23,6'd25,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd20,6'd22,6'd24,6'd31: Enemy_img = 4'd13;
//6'd19,6'd21,6'd23,6'd25,6'd27,6'd28,6'd29,6'd32,6'd34,6'd35,6'd39,6'd41,6'd43: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd30,6'd33: Enemy_img = 4'd9;
//6'd22,6'd24: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd27,6'd28,6'd35,6'd39,6'd41: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd30,6'd32,6'd33: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd10;
//6'd22,6'd24: Enemy_img = 4'd13;
//6'd20,6'd21,6'd23,6'd25,6'd26,6'd28,6'd35,6'd39,6'd41: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd30,6'd32,6'd33: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd10;
//6'd22,6'd24: Enemy_img = 4'd13;
//6'd21,6'd23,6'd25,6'd26,6'd28,6'd35,6'd39,6'd41: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd32: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd10;
//6'd24: Enemy_img = 4'd13;
//6'd22,6'd23,6'd25,6'd26,6'd28,6'd29,6'd34,6'd35,6'd39: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd24: Enemy_img = 4'd13;
//6'd23,6'd25,6'd26,6'd28,6'd29,6'd30,6'd33,6'd34,6'd39: Enemy_img = 4'd14;
//6'd35,6'd37,6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd31: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd28,6'd30,6'd32,6'd33: Enemy_img = 4'd14;
//6'd35,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd13;
//6'd32: Enemy_img = 4'd14;
//6'd25,6'd26,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd14;
//6'd26,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd37: Enemy_img = 4'd14;
//6'd27,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd36: Enemy_img = 4'd14;
//6'd28,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd13;
//6'd34,6'd39: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd13;
//6'd33,6'd39: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd36,6'd38,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd1;
//6'd38,6'd40: Enemy_img = 4'd14;
//6'd36,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd1;
//6'd28: Enemy_img = 4'd13;
//6'd36,6'd38,6'd40: Enemy_img = 4'd14;
//6'd35,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd1;
//6'd22,6'd28: Enemy_img = 4'd13;
//6'd21,6'd23,6'd29,6'd36,6'd39,6'd41: Enemy_img = 4'd14;
//6'd35,6'd37,6'd38,6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd1;
//6'd22,6'd28: Enemy_img = 4'd13;
//6'd17,6'd21,6'd29,6'd30,6'd31,6'd33,6'd37,6'd39,6'd41: Enemy_img = 4'd14;
//6'd34,6'd36,6'd38,6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd1;
//6'd23: Enemy_img = 4'd2;
//6'd29: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd28,6'd30,6'd31,6'd33,6'd37,6'd39: Enemy_img = 4'd14;
//6'd20,6'd34,6'd36,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd2;
//6'd18,6'd29: Enemy_img = 4'd13;
//6'd16,6'd17,6'd19,6'd20,6'd21,6'd26,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd40: Enemy_img = 4'd14;
//6'd35,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd24,6'd25: Enemy_img = 4'd2;
//6'd18,6'd20,6'd30: Enemy_img = 4'd13;
//6'd16,6'd17,6'd19,6'd21,6'd22,6'd23,6'd26,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd38,6'd40: Enemy_img = 4'd14;
//6'd35,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd25: Enemy_img = 4'd2;
//6'd18,6'd21,6'd23,6'd30: Enemy_img = 4'd13;
//6'd16,6'd17,6'd19,6'd20,6'd22,6'd24,6'd26,6'd27,6'd28,6'd29,6'd31,6'd34,6'd38,6'd39,6'd41: Enemy_img = 4'd14;
//6'd35,6'd37,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd25: Enemy_img = 4'd2;
//6'd32,6'd33: Enemy_img = 4'd9;
//6'd19,6'd21,6'd23: Enemy_img = 4'd13;
//6'd17,6'd18,6'd20,6'd22,6'd24,6'd26,6'd27,6'd28,6'd29,6'd35,6'd39: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd30,6'd32,6'd33: Enemy_img = 4'd9;
//6'd19,6'd21,6'd23,6'd24: Enemy_img = 4'd13;
//6'd17,6'd18,6'd20,6'd22,6'd25,6'd27,6'd28,6'd35,6'd39: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd2;
//6'd30,6'd32,6'd33: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd10;
//6'd20,6'd22,6'd24: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd21,6'd23,6'd25,6'd27,6'd28,6'd35,6'd36: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd1;
//6'd27: Enemy_img = 4'd2;
//6'd31: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd20,6'd22,6'd24: Enemy_img = 4'd13;
//6'd18,6'd19,6'd21,6'd23,6'd25,6'd26,6'd28,6'd29,6'd34,6'd35: Enemy_img = 4'd14;
//6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd2;
//6'd23,6'd25: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd24,6'd26,6'd27,6'd29,6'd30,6'd34,6'd35: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd2;
//6'd23,6'd25,6'd32,6'd33: Enemy_img = 4'd13;
//6'd21,6'd22,6'd24,6'd26,6'd27,6'd29,6'd30,6'd31,6'd34,6'd40: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd2;
//6'd26,6'd33: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd30,6'd40: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd2;
//6'd26: Enemy_img = 4'd13;
//6'd24,6'd25,6'd27,6'd28,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd14;
//6'd27,6'd28,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd14;
//6'd32,6'd33,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd35,6'd36: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd13;
//6'd33,6'd34,6'd36,6'd37: Enemy_img = 4'd14;
//6'd32,6'd35,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd1;
//6'd29,6'd34,6'd35,6'd37,6'd38: Enemy_img = 4'd14;
//6'd33,6'd36,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd1;
//6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd1;
//6'd34,6'd36,6'd37: Enemy_img = 4'd14;
//6'd32,6'd33,6'd35,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd1;
//6'd35,6'd37,6'd38: Enemy_img = 4'd14;
//6'd33,6'd34,6'd36,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd33: Enemy_img = 4'd1;
//6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//6'd31,6'd32,6'd34,6'd35,6'd37,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd1;
//6'd26: Enemy_img = 4'd13;
//6'd27,6'd31,6'd37,6'd39: Enemy_img = 4'd14;
//6'd28,6'd32,6'd33,6'd35,6'd36,6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd1;
//6'd26,6'd27: Enemy_img = 4'd13;
//6'd28,6'd29,6'd31,6'd32,6'd38: Enemy_img = 4'd14;
//6'd33,6'd34,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd1;
//6'd27,6'd28: Enemy_img = 4'd13;
//6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd39: Enemy_img = 4'd14;
//6'd34,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd1;
//6'd20,6'd28,6'd29: Enemy_img = 4'd13;
//6'd21,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd1;
//6'd24,6'd25: Enemy_img = 4'd2;
//6'd20,6'd29,6'd30: Enemy_img = 4'd13;
//6'd19,6'd28,6'd31,6'd35: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd1;
//6'd22,6'd23,6'd24: Enemy_img = 4'd2;
//6'd32,6'd33: Enemy_img = 4'd9;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd35,6'd36: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd1;
//6'd21,6'd24: Enemy_img = 4'd2;
//6'd33,6'd34: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd35,6'd36: Enemy_img = 4'd14;
//6'd37,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd2;
//6'd31,6'd34: Enemy_img = 4'd9;
//6'd32,6'd33: Enemy_img = 4'd10;
//6'd20: Enemy_img = 4'd13;
//6'd14,6'd16,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd36: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd2;
//6'd33: Enemy_img = 4'd10;
//6'd18,6'd20,6'd21,6'd23: Enemy_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd19,6'd22,6'd24,6'd25,6'd27,6'd28,6'd29,6'd35,6'd36: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd2;
//6'd18,6'd19,6'd21,6'd22,6'd24,6'd34,6'd35: Enemy_img = 4'd13;
//6'd15,6'd16,6'd17,6'd20,6'd23,6'd25,6'd26,6'd30,6'd31,6'd32,6'd36: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd2;
//6'd19,6'd20,6'd22,6'd23,6'd25,6'd35: Enemy_img = 4'd13;
//6'd16,6'd17,6'd18,6'd21,6'd24,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd2;
//6'd20,6'd21,6'd23,6'd24,6'd26: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd22,6'd25,6'd27,6'd28,6'd29,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd2;
//6'd21,6'd22,6'd24,6'd25,6'd27: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd23,6'd26,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd25,6'd26,6'd28: Enemy_img = 4'd13;
//6'd19,6'd20,6'd21,6'd23,6'd24,6'd27,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd27,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd33,6'd34: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd28,6'd29,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd1;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd33,6'd34: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd1;
//6'd25,6'd30,6'd31,6'd32,6'd35,6'd36: Enemy_img = 4'd14;
//6'd29,6'd33,6'd34,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd1;
//6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd30,6'd31,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd1;
//6'd35,6'd36: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd1;
//6'd28,6'd29,6'd37,6'd38: Enemy_img = 4'd14;
//6'd30,6'd31,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd1;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd41: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd1;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd41: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd9;
//6'd26,6'd27,6'd28: Enemy_img = 4'd13;
//6'd29,6'd30,6'd35,6'd36,6'd42: Enemy_img = 4'd14;
//6'd37,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd29,6'd30: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd36,6'd42: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd2;
//6'd34: Enemy_img = 4'd9;
//6'd32,6'd33: Enemy_img = 4'd10;
//6'd28,6'd29,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd2;
//6'd31,6'd32,6'd33: Enemy_img = 4'd9;
//6'd20: Enemy_img = 4'd13;
//6'd21,6'd26,6'd27,6'd28,6'd29,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd2;
//6'd21,6'd36: Enemy_img = 4'd13;
//6'd20,6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd26,6'd27: Enemy_img = 4'd2;
//6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd2;
//6'd24,6'd25: Enemy_img = 4'd13;
//6'd22,6'd23,6'd26,6'd27,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd2;
//6'd22,6'd26,6'd27: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd28,6'd29,6'd30: Enemy_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd35,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22,6'd25,6'd26,6'd27,6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd23,6'd24,6'd28,6'd29,6'd33,6'd34,6'd38,6'd39: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd28,6'd29: Enemy_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd36,6'd37: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd30: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd23,6'd24,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd26,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd22,6'd23: Enemy_img = 4'd13;
//6'd40: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd1;
//6'd22,6'd23,6'd41: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd1;
//6'd42: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd1;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd36,6'd37,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd27,6'd28,6'd29,6'd30,6'd36,6'd37: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd10;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38: Enemy_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd42: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd2;
//6'd22,6'd23,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd2;
//6'd22,6'd23: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40: Enemy_img = 4'd14;
//6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd13;
//6'd22,6'd23,6'd26,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd13;
//6'd23,6'd24,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_1 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd30: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd36,6'd37: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22,6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd38,6'd39: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19,6'd23,6'd24,6'd28,6'd29,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd1;
//6'd22,6'd26,6'd27: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd1;
//6'd24,6'd25,6'd33: Enemy_img = 4'd14;
//6'd22,6'd23,6'd26,6'd27,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd26,6'd27: Enemy_img = 4'd1;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd24,6'd25,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd1;
//6'd21: Enemy_img = 4'd13;
//6'd20,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd1;
//6'd31,6'd32,6'd33: Enemy_img = 4'd9;
//6'd20,6'd36,6'd37: Enemy_img = 4'd13;
//6'd21,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd1;
//6'd31,6'd32,6'd33: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd10;
//6'd36: Enemy_img = 4'd13;
//6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd9;
//6'd32,6'd33: Enemy_img = 4'd10;
//6'd27,6'd28,6'd29,6'd30,6'd36,6'd42: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd9;
//6'd29,6'd30: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd35,6'd36,6'd37,6'd42: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd2;
//6'd27,6'd28: Enemy_img = 4'd13;
//6'd25,6'd26,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd41: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd2;
//6'd24,6'd25,6'd26: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd41: Enemy_img = 4'd14;
//6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd2;
//6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd2;
//6'd37,6'd38: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd2;
//6'd35,6'd36: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd2;
//6'd32,6'd33,6'd34: Enemy_img = 4'd13;
//6'd30,6'd31,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd2;
//6'd30,6'd31,6'd32,6'd35,6'd36: Enemy_img = 4'd13;
//6'd25,6'd29,6'd33,6'd34,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd2;
//6'd25,6'd26,6'd33,6'd34: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd25,6'd26,6'd28,6'd29,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd33,6'd34: Enemy_img = 4'd13;
//6'd28,6'd30,6'd31,6'd32,6'd35: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd13;
//6'd27,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//2'd2: begin
//case(angle)
//// Enemy_type_2 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd9;
//6'd29,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd28,6'd31: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd9;
//6'd28,6'd31,6'd32: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd28,6'd32: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd6;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd9;
//6'd37: Enemy_img = 4'd11;
//6'd27,6'd33: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd9;
//6'd36,6'd37: Enemy_img = 4'd11;
//6'd27,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd6;
//6'd38: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd24,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd24,6'd25,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd10;
//6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd5;
//6'd28,6'd29: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd6;
//6'd28,6'd29: Enemy_img = 4'd10;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd10;
//6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd32,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd6;
//6'd38: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd6;
//6'd37: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd9;
//6'd26: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd9;
//6'd24,6'd26: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26: Enemy_img = 4'd9;
//6'd33: Enemy_img = 4'd11;
//6'd27,6'd28: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd6;
//6'd25,6'd26: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd11;
//6'd24,6'd27,6'd28: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd6;
//6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd9;
//6'd33,6'd35: Enemy_img = 4'd11;
//6'd24,6'd30,6'd31: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28: Enemy_img = 4'd9;
//6'd25,6'd29,6'd30: Enemy_img = 4'd14;
//6'd31,6'd32,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27: Enemy_img = 4'd9;
//6'd24,6'd28,6'd32,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd9;
//6'd24,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd29,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd27,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd22,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd10;
//6'd20,6'd21,6'd25,6'd26,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd23,6'd24,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd11;
//6'd20,6'd26,6'd31,6'd32: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd5;
//6'd28,6'd29,6'd30: Enemy_img = 4'd10;
//6'd19: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd38: Enemy_img = 4'd6;
//6'd29: Enemy_img = 4'd10;
//6'd39: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd6;
//6'd39: Enemy_img = 4'd11;
//6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd6;
//6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd28,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd35,6'd36,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd6;
//6'd43: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd5;
//6'd37: Enemy_img = 4'd6;
//6'd43: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd10;
//6'd42,6'd43: Enemy_img = 4'd14;
//6'd27,6'd29,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35: Enemy_img = 4'd10;
//6'd36: Enemy_img = 4'd11;
//6'd37,6'd38,6'd42: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd35: Enemy_img = 4'd11;
//6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd6;
//6'd35: Enemy_img = 4'd10;
//6'd24: Enemy_img = 4'd11;
//6'd32,6'd33,6'd37,6'd38: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd37,6'd40: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd9;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd41: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41: Enemy_img = 4'd9;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38: Enemy_img = 4'd14;
//6'd27,6'd28,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40: Enemy_img = 4'd9;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd9;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd42,6'd43: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd9;
//6'd26,6'd27,6'd28,6'd30,6'd31,6'd36,6'd37: Enemy_img = 4'd14;
//6'd32,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42: Enemy_img = 4'd9;
//6'd25,6'd26,6'd27,6'd37,6'd39,6'd40,6'd43: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd34,6'd36,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd6;
//6'd42,6'd43: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd11;
//6'd24,6'd25,6'd26,6'd41: Enemy_img = 4'd14;
//6'd28,6'd29,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34: Enemy_img = 4'd11;
//6'd23,6'd24,6'd25,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd11;
//6'd23,6'd24,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd14;
//6'd20,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd5;
//6'd34: Enemy_img = 4'd6;
//6'd40: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd10;
//6'd34: Enemy_img = 4'd11;
//6'd36,6'd37: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd35: Enemy_img = 4'd10;
//6'd34: Enemy_img = 4'd11;
//6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd25,6'd26,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd10;
//6'd32,6'd37,6'd39,6'd41: Enemy_img = 4'd14;
//6'd25,6'd26,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41: Enemy_img = 4'd9;
//6'd32,6'd33,6'd36,6'd38,6'd42: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd9;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd43: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd9;
//6'd23,6'd25: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd6;
//6'd39,6'd40,6'd43,6'd44: Enemy_img = 4'd9;
//6'd24: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd41,6'd42,6'd45: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd11;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd28,6'd29,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd45: Enemy_img = 4'd14;
//6'd29,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd38: Enemy_img = 4'd6;
//6'd37: Enemy_img = 4'd11;
//6'd29,6'd30: Enemy_img = 4'd14;
//6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd11;
//6'd29,6'd30: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd5;
//6'd32: Enemy_img = 4'd6;
//6'd29,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd9;
//6'd32: Enemy_img = 4'd10;
//6'd33: Enemy_img = 4'd11;
//6'd35,6'd36,6'd38,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd9;
//6'd31,6'd32,6'd34: Enemy_img = 4'd10;
//6'd33: Enemy_img = 4'd11;
//6'd36,6'd38,6'd45: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd9;
//6'd31,6'd34: Enemy_img = 4'd10;
//6'd36,6'd38,6'd46,6'd47: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd9;
//6'd32,6'd33,6'd35,6'd36,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd9;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd38,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd38,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd38,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd40: Enemy_img = 4'd6;
//6'd26,6'd39: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd30,6'd31,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd38: Enemy_img = 4'd6;
//6'd25,6'd26,6'd39,6'd40: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd30,6'd31,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd38: Enemy_img = 4'd11;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd14;
//6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd9;
//6'd36,6'd37,6'd39,6'd40,6'd42,6'd44: Enemy_img = 4'd14;
//6'd24,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd5;
//6'd29: Enemy_img = 4'd6;
//6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd9;
//6'd32,6'd33,6'd35,6'd38,6'd44: Enemy_img = 4'd14;
//6'd24: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd9;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd42,6'd43: Enemy_img = 4'd14;
//6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd9;
//6'd33,6'd34,6'd36,6'd40,6'd41: Enemy_img = 4'd14;
//6'd26,6'd27,6'd35,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd9;
//6'd30,6'd32: Enemy_img = 4'd10;
//6'd31: Enemy_img = 4'd11;
//6'd34,6'd36,6'd37,6'd40,6'd41: Enemy_img = 4'd14;
//6'd27,6'd28,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd9;
//6'd29,6'd30,6'd32: Enemy_img = 4'd10;
//6'd31: Enemy_img = 4'd11;
//6'd35,6'd38: Enemy_img = 4'd14;
//6'd24,6'd25,6'd27,6'd28,6'd36,6'd37,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd10;
//6'd32,6'd34,6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd27,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd39,6'd41: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd6;
//6'd40: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd11;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd19,6'd30,6'd31,6'd32,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd31,6'd32,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd28,6'd29: Enemy_img = 4'd6;
//6'd27: Enemy_img = 4'd11;
//6'd34,6'd35: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd11;
//6'd34,6'd35: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd9;
//6'd25,6'd26,6'd27,6'd28,6'd36,6'd38,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd9;
//6'd25,6'd28,6'd29,6'd35,6'd36,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd36,6'd37,6'd38: Enemy_img = 4'd9;
//6'd33,6'd35,6'd39: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd9;
//6'd32,6'd38: Enemy_img = 4'd14;
//6'd29,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd9;
//6'd30,6'd33,6'd38: Enemy_img = 4'd14;
//6'd21,6'd22,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd5;
//6'd35,6'd36,6'd37: Enemy_img = 4'd9;
//6'd29,6'd30,6'd31,6'd34: Enemy_img = 4'd14;
//6'd21,6'd33,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd5;
//6'd26: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd21,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd11;
//6'd33,6'd35,6'd37: Enemy_img = 4'd14;
//6'd21,6'd22,6'd34,6'd36,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd28,6'd31: Enemy_img = 4'd10;
//6'd29,6'd30: Enemy_img = 4'd11;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd10;
//6'd39,6'd40,6'd41: Enemy_img = 4'd11;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd6;
//6'd29: Enemy_img = 4'd10;
//6'd40: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd24,6'd27,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd6;
//6'd30: Enemy_img = 4'd11;
//6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32: Enemy_img = 4'd11;
//6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd11;
//6'd40,6'd41: Enemy_img = 4'd14;
//6'd20: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd9;
//6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd9;
//6'd32,6'd35: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd9;
//6'd31,6'd32,6'd35: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd30,6'd31,6'd35: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd22,6'd23,6'd24,6'd25,6'd30,6'd35: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd22,6'd29,6'd30,6'd35: Enemy_img = 4'd14;
//6'd26,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30,6'd36: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd11;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd5;
//6'd30: Enemy_img = 4'd10;
//6'd39: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd10;
//6'd28,6'd29: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd19,6'd20,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd10;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd19,6'd26,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd10;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd22,6'd23,6'd25,6'd26,6'd27,6'd31,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd11;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34: Enemy_img = 4'd11;
//6'd24,6'd25,6'd26,6'd27,6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd11;
//6'd20,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32: Enemy_img = 4'd11;
//6'd20,6'd21,6'd22,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd6;
//6'd21,6'd22: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd11;
//6'd23,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23: Enemy_img = 4'd9;
//6'd21,6'd24,6'd25,6'd27,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd26,6'd28,6'd30,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd9;
//6'd27,6'd28,6'd33,6'd34,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd29,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd9;
//6'd21,6'd22,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26: Enemy_img = 4'd9;
//6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd9;
//6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd27,6'd28,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd9;
//6'd23,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd26,6'd27,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd11;
//6'd24,6'd27,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd6;
//6'd29: Enemy_img = 4'd10;
//6'd40: Enemy_img = 4'd11;
//6'd26,6'd27,6'd31,6'd32: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd39,6'd40,6'd41: Enemy_img = 4'd11;
//6'd25,6'd26,6'd27: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31: Enemy_img = 4'd10;
//6'd28: Enemy_img = 4'd11;
//6'd22,6'd26,6'd27: Enemy_img = 4'd14;
//6'd23,6'd24,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd10;
//6'd21,6'd22: Enemy_img = 4'd14;
//6'd33,6'd35,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd5;
//6'd27: Enemy_img = 4'd6;
//6'd21: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27: Enemy_img = 4'd6;
//6'd21: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22: Enemy_img = 4'd14;
//6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd28,6'd29,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd11;
//6'd34,6'd35: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd28,6'd29: Enemy_img = 4'd6;
//6'd27: Enemy_img = 4'd11;
//6'd34,6'd35: Enemy_img = 4'd14;
//6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd19,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd11;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd27,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd6;
//6'd20,6'd21,6'd24,6'd25: Enemy_img = 4'd9;
//6'd40: Enemy_img = 4'd11;
//6'd19,6'd22,6'd23,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd27,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd20,6'd21,6'd22,6'd23,6'd24: Enemy_img = 4'd9;
//6'd39,6'd41: Enemy_img = 4'd11;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd27,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd22,6'd23,6'd24,6'd25: Enemy_img = 4'd9;
//6'd21,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd27,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25: Enemy_img = 4'd9;
//6'd22,6'd26,6'd28,6'd31,6'd32: Enemy_img = 4'd14;
//6'd27,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd10;
//6'd23,6'd25,6'd27,6'd32: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd31,6'd32: Enemy_img = 4'd10;
//6'd30: Enemy_img = 4'd11;
//6'd24,6'd25,6'd27,6'd28: Enemy_img = 4'd14;
//6'd35,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd10;
//6'd30: Enemy_img = 4'd11;
//6'd27,6'd28: Enemy_img = 4'd14;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27: Enemy_img = 4'd14;
//6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd5;
//6'd30: Enemy_img = 4'd6;
//6'd24: Enemy_img = 4'd14;
//6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//6'd32,6'd33,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd38: Enemy_img = 4'd11;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd38: Enemy_img = 4'd6;
//6'd25,6'd26,6'd39,6'd40: Enemy_img = 4'd11;
//6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd29,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd40: Enemy_img = 4'd6;
//6'd26,6'd39: Enemy_img = 4'd11;
//6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd29,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd27,6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd25,6'd27,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd23,6'd24,6'd27,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd9;
//6'd23,6'd24,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd21,6'd22,6'd27,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25: Enemy_img = 4'd9;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd26,6'd27,6'd29,6'd30,6'd32,6'd33: Enemy_img = 4'd14;
//6'd28,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd9;
//6'd31,6'd34: Enemy_img = 4'd10;
//6'd18,6'd19,6'd27,6'd29: Enemy_img = 4'd14;
//6'd28,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Enemy_img = 4'd9;
//6'd31,6'd33,6'd34: Enemy_img = 4'd10;
//6'd32: Enemy_img = 4'd11;
//6'd20,6'd27,6'd29: Enemy_img = 4'd14;
//6'd28,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd9;
//6'd33: Enemy_img = 4'd10;
//6'd32: Enemy_img = 4'd11;
//6'd22,6'd23,6'd24,6'd27,6'd29,6'd30: Enemy_img = 4'd14;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd14;
//6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd5;
//6'd33: Enemy_img = 4'd6;
//6'd29,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30: Enemy_img = 4'd14;
//6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd11;
//6'd29,6'd30: Enemy_img = 4'd14;
//6'd26: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd38: Enemy_img = 4'd6;
//6'd37: Enemy_img = 4'd11;
//6'd29,6'd30: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd27,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd27,6'd28,6'd32,6'd33,6'd34,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd6;
//6'd24: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd27,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd6;
//6'd23,6'd25: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd6;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd26,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd26,6'd27,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd10;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd32: Enemy_img = 4'd14;
//6'd27,6'd37,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd9;
//6'd32,6'd34,6'd35: Enemy_img = 4'd10;
//6'd33: Enemy_img = 4'd11;
//6'd26,6'd29: Enemy_img = 4'd14;
//6'd23,6'd24,6'd27,6'd28,6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd9;
//6'd32,6'd34: Enemy_img = 4'd10;
//6'd33: Enemy_img = 4'd11;
//6'd23,6'd24,6'd27,6'd28,6'd30: Enemy_img = 4'd14;
//6'd29,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27: Enemy_img = 4'd9;
//6'd23,6'd24,6'd28,6'd30,6'd31: Enemy_img = 4'd14;
//6'd22,6'd29,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd9;
//6'd21,6'd22,6'd28,6'd29,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd5;
//6'd35: Enemy_img = 4'd6;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28: Enemy_img = 4'd9;
//6'd20,6'd26,6'd29,6'd31,6'd32: Enemy_img = 4'd14;
//6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23: Enemy_img = 4'd9;
//6'd20,6'd22,6'd24,6'd25,6'd27,6'd28: Enemy_img = 4'd14;
//6'd31,6'd32,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd11;
//6'd23,6'd24: Enemy_img = 4'd14;
//6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34: Enemy_img = 4'd11;
//6'd23,6'd24,6'd25: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd6;
//6'd34: Enemy_img = 4'd11;
//6'd24,6'd25,6'd26: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27: Enemy_img = 4'd14;
//6'd37,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28: Enemy_img = 4'd14;
//6'd30,6'd31,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//6'd24,6'd25,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//6'd25,6'd26,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd26,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd26,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd27,6'd37,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd6;
//6'd35: Enemy_img = 4'd10;
//6'd24: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd10;
//6'd23,6'd24,6'd25: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd26,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24: Enemy_img = 4'd6;
//6'd33,6'd35,6'd36: Enemy_img = 4'd10;
//6'd34: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd27,6'd37,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd11;
//6'd27,6'd29,6'd31: Enemy_img = 4'd14;
//6'd26,6'd28,6'd30,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38: Enemy_img = 4'd6;
//6'd26,6'd27,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd30,6'd31,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd5;
//6'd27,6'd28,6'd29: Enemy_img = 4'd9;
//6'd30,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd25,6'd26,6'd31,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Enemy_img = 4'd9;
//6'd26,6'd31,6'd34: Enemy_img = 4'd14;
//6'd25,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd9;
//6'd26,6'd32: Enemy_img = 4'd14;
//6'd25,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd30: Enemy_img = 4'd9;
//6'd25,6'd29,6'd31: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27: Enemy_img = 4'd9;
//6'd24,6'd28,6'd29,6'd35,6'd36,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25: Enemy_img = 4'd9;
//6'd24,6'd26,6'd28,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31: Enemy_img = 4'd11;
//6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd6;
//6'd30: Enemy_img = 4'd11;
//6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd6;
//6'd29,6'd31: Enemy_img = 4'd11;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22: Enemy_img = 4'd14;
//6'd32,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd23,6'd24,6'd33,6'd37,6'd38,6'd39,6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd10;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd25,6'd26,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd10;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd26,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd6;
//6'd34: Enemy_img = 4'd10;
//6'd35,6'd36: Enemy_img = 4'd11;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//6'd27,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd5;
//6'd26: Enemy_img = 4'd6;
//6'd35: Enemy_img = 4'd10;
//6'd25: Enemy_img = 4'd11;
//6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd6;
//6'd25: Enemy_img = 4'd11;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd11;
//6'd28,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd37: Enemy_img = 4'd14;
//6'd28,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd32,6'd33: Enemy_img = 4'd9;
//6'd29,6'd31,6'd34,6'd35,6'd43: Enemy_img = 4'd14;
//6'd28,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd9;
//6'd29,6'd35,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33: Enemy_img = 4'd9;
//6'd29,6'd30,6'd34,6'd41: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd9;
//6'd29,6'd30,6'd33: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd9;
//6'd29,6'd32: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd9;
//6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd6;
//6'd28: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd11;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd6;
//6'd27: Enemy_img = 4'd11;
//6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd10;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd6;
//6'd36,6'd37: Enemy_img = 4'd10;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd5;
//6'd36,6'd37: Enemy_img = 4'd11;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd10;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd45: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd44,6'd45: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd6;
//6'd27: Enemy_img = 4'd11;
//6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd9;
//6'd28,6'd29: Enemy_img = 4'd11;
//6'd31,6'd32,6'd33,6'd34,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd9;
//6'd28: Enemy_img = 4'd11;
//6'd32,6'd38: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36: Enemy_img = 4'd9;
//6'd33,6'd37: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd9;
//6'd33,6'd34,6'd37: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd9;
//6'd34,6'd37: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd9;
//6'd34: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd9;
//6'd34,6'd36: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_2 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd11;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26: Enemy_img = 4'd6;
//6'd25: Enemy_img = 4'd11;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd39: Enemy_img = 4'd6;
//6'd35: Enemy_img = 4'd10;
//6'd25: Enemy_img = 4'd11;
//6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd5;
//6'd34,6'd35,6'd36: Enemy_img = 4'd10;
//6'd45: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd11;
//6'd32,6'd33,6'd38,6'd44: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd10;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd43,6'd44: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd40,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39: Enemy_img = 4'd14;
//6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd9;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd40: Enemy_img = 4'd14;
//6'd28,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd9;
//6'd20,6'd21,6'd22,6'd32,6'd36,6'd40: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38: Enemy_img = 4'd9;
//6'd34,6'd35,6'd39: Enemy_img = 4'd14;
//6'd25,6'd32,6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30: Enemy_img = 4'd6;
//6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd9;
//6'd29,6'd31: Enemy_img = 4'd11;
//6'd33,6'd34,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32: Enemy_img = 4'd6;
//6'd38,6'd39: Enemy_img = 4'd9;
//6'd30: Enemy_img = 4'd11;
//6'd36,6'd37,6'd40: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40: Enemy_img = 4'd9;
//6'd31: Enemy_img = 4'd11;
//6'd36,6'd37: Enemy_img = 4'd14;
//6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd9;
//6'd38,6'd40: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd9;
//6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//2'd3: begin
//case(angle)
//// Enemy_type_3 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd50,6'd51,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd13;
//6'd26,6'd27,6'd29,6'd30,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69: Enemy_img = 4'd14;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29: Enemy_img = 4'd13;
//6'd25,6'd26,6'd30,6'd31,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd61,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd13;
//6'd25,6'd26,6'd30,6'd31,6'd32,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd60,6'd62,6'd70: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd31,6'd32,6'd33,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd43,6'd59,6'd63,6'd69: Enemy_img = 4'd13;
//6'd24,6'd25,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd32,6'd42,6'd44,6'd58,6'd63,6'd69: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd31,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd32,6'd33,6'd35,6'd36,6'd41,6'd45,6'd56,6'd57,6'd60,6'd61,6'd64: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38,6'd39,6'd40,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd62,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd43,6'd52,6'd54,6'd55,6'd59,6'd60,6'd61,6'd64,6'd68: Enemy_img = 4'd13;
//6'd23,6'd24,6'd28,6'd35,6'd39,6'd40,6'd42,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd58,6'd62,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd29,6'd30,6'd34,6'd36,6'd37,6'd40,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd67: Enemy_img = 4'd13;
//6'd23,6'd24,6'd28,6'd31,6'd32,6'd35,6'd38,6'd39,6'd42,6'd45,6'd56,6'd57,6'd63,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd32,6'd34,6'd35,6'd36,6'd37,6'd39,6'd42,6'd43,6'd44,6'd45,6'd56,6'd62,6'd65,6'd67: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd31,6'd38,6'd41,6'd46,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd39,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63: Enemy_img = 4'd13;
//6'd22,6'd23,6'd31,6'd37,6'd38,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd51,6'd58,6'd61,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd41,6'd42,6'd44,6'd45,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57,6'd66: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd43,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd52,6'd53,6'd58,6'd59: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd38,6'd42,6'd61,6'd62,6'd63,6'd64,6'd67: Enemy_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd36,6'd37,6'd40,6'd41,6'd43,6'd44,6'd49,6'd50,6'd55,6'd56,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd51,6'd52,6'd57,6'd58: Enemy_img = 4'd9;
//6'd32,6'd37,6'd40,6'd42,6'd43,6'd48,6'd49,6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd39,6'd41,6'd65,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd52,6'd58: Enemy_img = 4'd9;
//6'd45,6'd51,6'd57: Enemy_img = 4'd10;
//6'd40,6'd42,6'd43,6'd48,6'd49,6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68: Enemy_img = 4'd13;
//6'd39,6'd41,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//endcase
//end
//6'd62: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd38,6'd44,6'd47,6'd50,6'd53,6'd56,6'd59,6'd68,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd45,6'd46,6'd51,6'd52,6'd57,6'd58: Enemy_img = 4'd10;
//default: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//endcase
//end
//6'd63: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd38,6'd44,6'd47,6'd50,6'd53,6'd56,6'd59,6'd68,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd46,6'd52,6'd58: Enemy_img = 4'd9;
//6'd45,6'd51,6'd57: Enemy_img = 4'd10;
//6'd48,6'd54,6'd60: Enemy_img = 4'd13;
//default: Enemy_img = 4'd14;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd51,6'd52,6'd57,6'd58: Enemy_img = 4'd9;
//6'd48,6'd54,6'd60: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd51,6'd57: Enemy_img = 4'd9;
//6'd48,6'd54,6'd60: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd22,6'd46,6'd52,6'd58,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd55,6'd61: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50,6'd56,6'd62,6'd63,6'd64,6'd65,6'd67,6'd69: Enemy_img = 4'd14;
//6'd20,6'd21,6'd38,6'd46,6'd47,6'd52,6'd53,6'd58,6'd59,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd55,6'd61: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd50,6'd51,6'd56,6'd57,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//6'd21,6'd38,6'd68,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd22,6'd39,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd22,6'd39,6'd65,6'd68,6'd69,6'd70,6'd72,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68,6'd69,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd23,6'd40,6'd47,6'd48,6'd49,6'd50,6'd51,6'd65,6'd70,6'd72,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd68,6'd73,6'd74: Enemy_img = 4'd14;
//6'd23,6'd40,6'd46,6'd52,6'd53,6'd54,6'd55,6'd64,6'd66,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd65,6'd68,6'd69,6'd70,6'd71,6'd73: Enemy_img = 4'd14;
//6'd23,6'd40,6'd41,6'd45,6'd52,6'd56,6'd57,6'd64,6'd66,6'd72,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd41,6'd45,6'd46,6'd47,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd24,6'd39,6'd40,6'd42,6'd44,6'd48,6'd49,6'd50,6'd51,6'd52,6'd58,6'd63,6'd67,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd24,6'd34,6'd39,6'd43,6'd48,6'd59,6'd63,6'd67,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd24,6'd33,6'd48,6'd60,6'd62,6'd68,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd43,6'd44,6'd45,6'd46,6'd47,6'd56,6'd57,6'd58,6'd59,6'd60,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd25,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd49,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd67: Enemy_img = 4'd14;
//6'd25,6'd31,6'd45,6'd46,6'd47,6'd48,6'd50,6'd55,6'd61,6'd66,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd25,6'd31,6'd50,6'd55,6'd58,6'd59,6'd60,6'd61,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd26,6'd30,6'd50,6'd55,6'd58,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//6'd26,6'd30,6'd50,6'd55,6'd58,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd64: Enemy_img = 4'd14;
//6'd27,6'd29,6'd50,6'd55,6'd58,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd52,6'd53,6'd54,6'd62,6'd63: Enemy_img = 4'd14;
//6'd27,6'd29,6'd55,6'd56,6'd57,6'd60,6'd61,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd28,6'd50,6'd51,6'd58,6'd59,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd58,6'd60,6'd61: Enemy_img = 4'd14;
//6'd28,6'd52,6'd53,6'd56,6'd57,6'd59,6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd56,6'd57,6'd58: Enemy_img = 4'd14;
//6'd54,6'd55,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd14;
//6'd54,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd57,6'd58,6'd59: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd60,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd57,6'd58,6'd59: Enemy_img = 4'd14;
//6'd56,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd57,6'd58: Enemy_img = 4'd14;
//6'd56,6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56: Enemy_img = 4'd14;
//6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56: Enemy_img = 4'd14;
//6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd70,6'd71: Enemy_img = 4'd14;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd99,6'd100,6'd101: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd61,6'd62,6'd68,6'd69,6'd70,6'd71,6'd72,6'd96,6'd102: Enemy_img = 4'd14;
//6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd97,6'd98: Enemy_img = 4'd13;
//6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd64,6'd65,6'd66,6'd69,6'd70,6'd94,6'd95,6'd96,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd94,6'd95,6'd96: Enemy_img = 4'd13;
//6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd89,6'd90,6'd91,6'd92,6'd93,6'd97,6'd98: Enemy_img = 4'd14;
//6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd92,6'd93: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd64,6'd89,6'd90,6'd91: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86,6'd87,6'd88,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd57,6'd58,6'd87,6'd88: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd58,6'd59,6'd64,6'd84,6'd85,6'd86: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd63,6'd82,6'd83,6'd84: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd57,6'd61,6'd63,6'd80,6'd81: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd58,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd56,6'd57,6'd58,6'd62,6'd77,6'd78,6'd79: Enemy_img = 4'd13;
//6'd22,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd59,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd56,6'd57,6'd58,6'd59,6'd75,6'd76,6'd77: Enemy_img = 4'd13;
//6'd22,6'd23,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd55,6'd56,6'd59,6'd60,6'd64,6'd73,6'd74: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd57,6'd58,6'd61,6'd62,6'd65,6'd66,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd51,6'd57,6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd49,6'd53,6'd54,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68,6'd69: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd55,6'd56,6'd59,6'd64,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd42,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd13;
//6'd22,6'd23,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd50,6'd51,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd9;
//6'd24,6'd25,6'd39,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd13;
//6'd22,6'd23,6'd26,6'd27,6'd28,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd49,6'd50,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd73,6'd74,6'd75,6'd76,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd41,6'd42,6'd50,6'd59,6'd60: Enemy_img = 4'd13;
//6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd43,6'd44,6'd47,6'd48,6'd49,6'd54,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd71,6'd72,6'd76,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd9;
//6'd56,6'd57,6'd58: Enemy_img = 4'd10;
//6'd24,6'd25,6'd26,6'd27,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd54,6'd60: Enemy_img = 4'd13;
//6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd45,6'd46,6'd61,6'd62,6'd63,6'd64,6'd65,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77: Enemy_img = 4'd14;
//6'd68,6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd9;
//6'd57,6'd58: Enemy_img = 4'd10;
//6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44,6'd45,6'd54,6'd55,6'd60: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd29,6'd37,6'd38,6'd40,6'd48,6'd49,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd69,6'd73,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd58: Enemy_img = 4'd9;
//6'd51,6'd52,6'd57: Enemy_img = 4'd10;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd35,6'd36,6'd38,6'd44,6'd48,6'd49,6'd54,6'd61: Enemy_img = 4'd13;
//6'd22,6'd23,6'd29,6'd34,6'd37,6'd40,6'd41,6'd42,6'd43,6'd55,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd69,6'd70,6'd73,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd58: Enemy_img = 4'd9;
//6'd51,6'd52: Enemy_img = 4'd10;
//6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd41,6'd42,6'd48,6'd49,6'd54,6'd55,6'd62: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd34,6'd37,6'd40,6'd43,6'd44,6'd56,6'd63,6'd64,6'd65,6'd68,6'd69,6'd73,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd59,6'd70,6'd71,6'd72,6'd74,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd52,6'd53: Enemy_img = 4'd9;
//6'd25,6'd26,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd38,6'd42,6'd43,6'd48,6'd49,6'd55,6'd62,6'd80,6'd81: Enemy_img = 4'd13;
//6'd23,6'd24,6'd27,6'd31,6'd37,6'd40,6'd41,6'd50,6'd56,6'd63,6'd64,6'd65,6'd69,6'd70,6'd71,6'd75,6'd79,6'd82: Enemy_img = 4'd14;
//6'd59,6'd60,6'd67,6'd72,6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53: Enemy_img = 4'd9;
//6'd46,6'd47: Enemy_img = 4'd10;
//6'd25,6'd26,6'd29,6'd33,6'd34,6'd38,6'd42,6'd43,6'd44,6'd49,6'd56,6'd78,6'd79: Enemy_img = 4'd13;
//6'd23,6'd24,6'd27,6'd28,6'd30,6'd31,6'd35,6'd36,6'd37,6'd40,6'd41,6'd50,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd70,6'd71,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd67,6'd68,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd53: Enemy_img = 4'd9;
//6'd46: Enemy_img = 4'd10;
//6'd25,6'd26,6'd27,6'd30,6'd38,6'd41,6'd49,6'd57: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd28,6'd29,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd42,6'd43,6'd44,6'd50,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd71,6'd72,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd54,6'd55,6'd67,6'd69,6'd75,6'd76,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd9;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd50: Enemy_img = 4'd13;
//6'd23,6'd24,6'd31,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd51,6'd52,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd67,6'd70,6'd75,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd9;
//6'd25,6'd26,6'd27,6'd31,6'd33,6'd51: Enemy_img = 4'd13;
//6'd23,6'd24,6'd28,6'd29,6'd30,6'd34,6'd35,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd73,6'd77: Enemy_img = 4'd14;
//6'd48,6'd49,6'd67,6'd71,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd29,6'd30,6'd36,6'd37,6'd38: Enemy_img = 4'd13;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd31,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd67,6'd72,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd34,6'd35,6'd36: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd29,6'd30,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd72,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd63,6'd64,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd32,6'd33,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd41,6'd51,6'd52,6'd56,6'd65,6'd66,6'd67,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd42,6'd55,6'd56,6'd66,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd27,6'd28,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd46,6'd47,6'd48,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd43,6'd44,6'd50,6'd53,6'd54,6'd66,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd48,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd62,6'd63,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd44,6'd45,6'd49,6'd53,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50,6'd51,6'd52,6'd55,6'd58,6'd59,6'd60,6'd62,6'd63,6'd65,6'd66,6'd67,6'd70: Enemy_img = 4'd14;
//6'd45,6'd46,6'd49,6'd53,6'd54,6'd56,6'd57,6'd61,6'd64,6'd69,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd66,6'd70: Enemy_img = 4'd14;
//6'd26,6'd45,6'd48,6'd49,6'd54,6'd55,6'd56,6'd61,6'd62,6'd65,6'd68,6'd69,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd69,6'd70: Enemy_img = 4'd14;
//6'd25,6'd26,6'd45,6'd53,6'd54,6'd56,6'd57,6'd62,6'd65,6'd68,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd68,6'd69: Enemy_img = 4'd14;
//6'd25,6'd26,6'd45,6'd52,6'd53,6'd57,6'd62,6'd63,6'd64,6'd67,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd68: Enemy_img = 4'd14;
//6'd27,6'd28,6'd57,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66: Enemy_img = 4'd14;
//6'd28,6'd29,6'd40,6'd58,6'd65,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd29,6'd40,6'd64,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd30,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd31,6'd39,6'd63,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd61,6'd62,6'd63,6'd67,6'd68: Enemy_img = 4'd14;
//6'd32,6'd39,6'd64,6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68: Enemy_img = 4'd14;
//6'd33,6'd39,6'd66,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd33,6'd39,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd34,6'd35,6'd39,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd67,6'd68: Enemy_img = 4'd14;
//6'd37,6'd39,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd14;
//6'd38,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd14;
//6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd74,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd75,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd75,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd75,6'd87,6'd88,6'd89,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd76,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd92: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92: Enemy_img = 4'd13;
//6'd45,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd96: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91: Enemy_img = 4'd13;
//6'd46,6'd47,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd74,6'd75,6'd76,6'd77,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89,6'd93: Enemy_img = 4'd13;
//6'd47,6'd48,6'd51,6'd52,6'd53,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd85,6'd88,6'd92,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd46,6'd49,6'd50,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd92,6'd93: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd87,6'd91,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd91,6'd92,6'd94,6'd95: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51,6'd54,6'd55,6'd56,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd86,6'd90,6'd93,6'd96,6'd97: Enemy_img = 4'd14;
//6'd47,6'd50,6'd52,6'd53,6'd57,6'd58,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd90,6'd91,6'd93,6'd94,6'd95: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd89,6'd92,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd65,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd58,6'd59,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd71,6'd78,6'd79,6'd80,6'd81,6'd84,6'd91,6'd97,6'd98: Enemy_img = 4'd14;
//6'd47,6'd60,6'd61,6'd64,6'd65,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd87,6'd91,6'd94,6'd95,6'd96: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd80,6'd83,6'd90,6'd92,6'd93,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd47,6'd48,6'd53,6'd61,6'd62,6'd64,6'd65,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd87,6'd95,6'd96: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd59,6'd60,6'd61,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82,6'd86,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd48,6'd53,6'd55,6'd56,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd86,6'd87,6'd92,6'd93,6'd97,6'd98: Enemy_img = 4'd13;
//6'd49,6'd52,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd85,6'd88,6'd90,6'd91,6'd94,6'd95,6'd96,6'd99,6'd100: Enemy_img = 4'd14;
//6'd48,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd62,6'd63,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd88,6'd92,6'd93,6'd96,6'd97,6'd98: Enemy_img = 4'd13;
//6'd55,6'd56,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd84,6'd85,6'd87,6'd90,6'd91,6'd94,6'd95,6'd99,6'd100: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd57,6'd58,6'd62,6'd66,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd88,6'd89,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd13;
//6'd50,6'd51,6'd56,6'd57,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd93,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd49,6'd52,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd65,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd13;
//6'd50,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd71,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd85,6'd86,6'd93,6'd94,6'd100,6'd101: Enemy_img = 4'd14;
//6'd49,6'd51,6'd55,6'd56,6'd59,6'd60,6'd64,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd9;
//6'd84,6'd86,6'd87,6'd88,6'd97,6'd98,6'd99: Enemy_img = 4'd13;
//6'd50,6'd53,6'd54,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd70,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd89,6'd92,6'd93,6'd94,6'd95,6'd96,6'd100,6'd101: Enemy_img = 4'd14;
//6'd48,6'd49,6'd51,6'd55,6'd56,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd9;
//6'd76: Enemy_img = 4'd10;
//6'd70,6'd78,6'd79,6'd80,6'd84,6'd87,6'd88,6'd89,6'd90,6'd100: Enemy_img = 4'd13;
//6'd50,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd69,6'd81,6'd82,6'd83,6'd85,6'd86,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd101,6'd102: Enemy_img = 4'd14;
//6'd48,6'd49,6'd51,6'd55,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd9;
//6'd76,6'd77: Enemy_img = 4'd10;
//6'd71,6'd72,6'd73,6'd80,6'd81,6'd82,6'd85,6'd87,6'd88: Enemy_img = 4'd13;
//6'd50,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd66,6'd67,6'd68,6'd69,6'd70,6'd83,6'd86,6'd89,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd49,6'd54,6'd55,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78: Enemy_img = 4'd9;
//6'd76: Enemy_img = 4'd10;
//6'd73,6'd74,6'd85: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd65,6'd66,6'd67,6'd72,6'd80,6'd81,6'd82,6'd83,6'd86,6'd87,6'd88,6'd89,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd77,6'd78: Enemy_img = 4'd9;
//6'd74,6'd75,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd13;
//6'd52,6'd53,6'd63,6'd64,6'd65,6'd66,6'd73,6'd84,6'd86,6'd87,6'd88,6'd89,6'd102,6'd103: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd54,6'd55,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd77: Enemy_img = 4'd9;
//6'd72: Enemy_img = 4'd10;
//6'd66,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd13;
//6'd52,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd84,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd49,6'd53,6'd54,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd9;
//6'd72,6'd73: Enemy_img = 4'd10;
//6'd66,6'd67,6'd68,6'd75,6'd79,6'd80,6'd81,6'd82,6'd83,6'd86: Enemy_img = 4'd13;
//6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd84,6'd87,6'd88: Enemy_img = 4'd14;
//6'd49,6'd51,6'd52,6'd53,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd9;
//6'd72: Enemy_img = 4'd10;
//6'd69: Enemy_img = 4'd13;
//6'd51,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd76,6'd78,6'd79,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd48,6'd49,6'd52,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd73,6'd74: Enemy_img = 4'd9;
//6'd70,6'd76,6'd80,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd68,6'd69,6'd77,6'd81,6'd82,6'd87: Enemy_img = 4'd14;
//6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd73: Enemy_img = 4'd9;
//6'd70,6'd71,6'd75,6'd79: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd69,6'd76,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd47,6'd51,6'd52,6'd53,6'd57,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66: Enemy_img = 4'd9;
//6'd67,6'd68: Enemy_img = 4'd10;
//6'd62,6'd63,6'd71,6'd75,6'd78: Enemy_img = 4'd13;
//6'd50,6'd51,6'd59,6'd60,6'd61,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd49,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd9;
//6'd67,6'd68: Enemy_img = 4'd10;
//6'd64,6'd65,6'd73,6'd74,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd71,6'd72,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd57,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69: Enemy_img = 4'd9;
//6'd65,6'd66,6'd72,6'd73,6'd77: Enemy_img = 4'd13;
//6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd71,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd9;
//6'd66,6'd67,6'd71,6'd72,6'd73: Enemy_img = 4'd13;
//6'd46,6'd47,6'd51,6'd52,6'd54,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd49,6'd50,6'd53,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd65,6'd66,6'd67,6'd73,6'd75: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd50,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd71,6'd72,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd64,6'd65,6'd66,6'd67,6'd70,6'd75: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd68,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd42,6'd48,6'd49,6'd52,6'd57,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd63,6'd64,6'd65,6'd66,6'd72,6'd75: Enemy_img = 4'd13;
//6'd43,6'd44,6'd47,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd49,6'd52,6'd53,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd65,6'd68,6'd71,6'd72,6'd74: Enemy_img = 4'd13;
//6'd46,6'd50,6'd51,6'd54,6'd58,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd47,6'd49,6'd52,6'd53,6'd55,6'd56,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd45,6'd50,6'd51,6'd53,6'd57,6'd58,6'd59,6'd65,6'd66,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd52,6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd64,6'd71,6'd72: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52,6'd56,6'd57,6'd58,6'd68,6'd69,6'd70,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd14;
//6'd46,6'd48,6'd51,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd67: Enemy_img = 4'd13;
//6'd49,6'd50,6'd55,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd14;
//6'd48,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd13;
//6'd49,6'd50,6'd54,6'd55,6'd56,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd14;
//6'd47,6'd48,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd66,6'd72,6'd73,6'd74: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd66: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd67: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd67: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd70,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd61,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd65: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd62,6'd63,6'd64,6'd66,6'd67,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd43,6'd58,6'd59,6'd60,6'd61,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd64: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd52,6'd61,6'd62,6'd63,6'd65,6'd66,6'd91,6'd92: Enemy_img = 4'd14;
//6'd42,6'd59,6'd60,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd63: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd60,6'd61,6'd62,6'd64,6'd65: Enemy_img = 4'd14;
//6'd41,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd62,6'd63: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd61,6'd64: Enemy_img = 4'd14;
//6'd40,6'd65,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd62: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd63: Enemy_img = 4'd14;
//6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd43,6'd44,6'd45: Enemy_img = 4'd14;
//6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd14;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd40,6'd41: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd13;
//6'd36,6'd37,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd13;
//6'd36,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd13;
//6'd35: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd13;
//6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd83: Enemy_img = 4'd14;
//6'd59,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd82,6'd83: Enemy_img = 4'd14;
//6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd13;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd79: Enemy_img = 4'd13;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd81: Enemy_img = 4'd13;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd81,6'd83: Enemy_img = 4'd13;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd80,6'd82,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd80,6'd83,6'd84,6'd85: Enemy_img = 4'd13;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd79,6'd81,6'd82,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd13;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd79,6'd81,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd13;
//6'd75,6'd78,6'd79,6'd81,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd79,6'd81,6'd88: Enemy_img = 4'd13;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd81,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd13;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd80,6'd82,6'd85,6'd86,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd77,6'd78,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd13;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd80,6'd81,6'd82,6'd85,6'd92,6'd93: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd78,6'd80,6'd83,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd13;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd77,6'd79,6'd82,6'd84,6'd85,6'd93,6'd94: Enemy_img = 4'd14;
//6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd78,6'd80,6'd83,6'd84: Enemy_img = 4'd13;
//6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd77,6'd79,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd13;
//6'd60,6'd61,6'd62,6'd73,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd13;
//6'd59,6'd60,6'd70,6'd71,6'd76,6'd77,6'd78,6'd81,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd13;
//6'd58,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd78: Enemy_img = 4'd14;
//6'd57,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd80,6'd81,6'd82: Enemy_img = 4'd13;
//6'd55,6'd56,6'd58,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd78,6'd79,6'd83: Enemy_img = 4'd14;
//6'd57,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd78,6'd80,6'd81: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd79,6'd82,6'd83: Enemy_img = 4'd14;
//6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd79: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd49,6'd50,6'd56,6'd57,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74,6'd75,6'd76,6'd79: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd55,6'd56,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd71,6'd72,6'd77,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd42,6'd48,6'd49,6'd53,6'd54,6'd57,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69: Enemy_img = 4'd9;
//6'd70: Enemy_img = 4'd10;
//6'd73,6'd74,6'd77: Enemy_img = 4'd13;
//6'd39,6'd43,6'd44,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd60,6'd61,6'd62,6'd64,6'd65,6'd75,6'd76,6'd78,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd55,6'd56,6'd59,6'd63,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69: Enemy_img = 4'd9;
//6'd70,6'd71,6'd72: Enemy_img = 4'd10;
//6'd77,6'd78,6'd81: Enemy_img = 4'd13;
//6'd39,6'd45,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd61,6'd64,6'd74,6'd75,6'd76,6'd79,6'd82,6'd83: Enemy_img = 4'd14;
//6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd56,6'd59,6'd62,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73: Enemy_img = 4'd9;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd81: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd60,6'd61,6'd64,6'd80,6'd82,6'd83: Enemy_img = 4'd14;
//6'd39,6'd40,6'd46,6'd55,6'd59,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd9;
//6'd65,6'd66,6'd68,6'd69,6'd75,6'd76,6'd77,6'd81: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd56,6'd57,6'd60,6'd63,6'd64,6'd67,6'd82,6'd83: Enemy_img = 4'd14;
//6'd40,6'd49,6'd50,6'd51,6'd55,6'd58,6'd59,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd9;
//6'd70,6'd71,6'd79: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd56,6'd57,6'd58,6'd63,6'd64,6'd65,6'd68,6'd69,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd40,6'd41,6'd48,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66: Enemy_img = 4'd9;
//6'd70,6'd71,6'd77: Enemy_img = 4'd13;
//6'd43,6'd44,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd62,6'd63,6'd72,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd41,6'd42,6'd45,6'd46,6'd47,6'd49,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67: Enemy_img = 4'd9;
//6'd68,6'd69: Enemy_img = 4'd10;
//6'd73,6'd76: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd72,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd59,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd70: Enemy_img = 4'd9;
//6'd68,6'd69: Enemy_img = 4'd10;
//6'd72,6'd76: Enemy_img = 4'd13;
//6'd45,6'd46,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd43,6'd44,6'd47,6'd51,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65,6'd66,6'd72,6'd75: Enemy_img = 4'd13;
//6'd45,6'd46,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd44,6'd47,6'd51,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71: Enemy_img = 4'd9;
//6'd67,6'd68,6'd75: Enemy_img = 4'd13;
//6'd46,6'd49,6'd52,6'd53,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd44,6'd45,6'd47,6'd50,6'd51,6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd72,6'd75: Enemy_img = 4'd13;
//6'd46,6'd49,6'd50,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd66,6'd67,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd44,6'd45,6'd47,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65: Enemy_img = 4'd9;
//6'd69,6'd71,6'd72: Enemy_img = 4'd13;
//6'd46,6'd49,6'd50,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd70,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd45,6'd47,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65: Enemy_img = 4'd9;
//6'd66,6'd67: Enemy_img = 4'd10;
//6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd51,6'd53,6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd9;
//6'd66: Enemy_img = 4'd10;
//6'd60,6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52,6'd56,6'd57,6'd58,6'd59,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd14;
//6'd46,6'd47,6'd51,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd9;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd75: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd50,6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd9;
//6'd65,6'd66,6'd72,6'd75: Enemy_img = 4'd13;
//6'd49,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd70,6'd71,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd46,6'd47,6'd50,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd70,6'd72,6'd75: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd71,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd47,6'd54,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd71,6'd72,6'd73,6'd75: Enemy_img = 4'd13;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd70,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd47,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd76: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd61,6'd62,6'd63,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd13;
//6'd47,6'd56,6'd57,6'd58,6'd62,6'd63,6'd76,6'd77,6'd78,6'd79,6'd80,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd65,6'd66,6'd70: Enemy_img = 4'd13;
//6'd47,6'd48,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd67,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd50,6'd51,6'd52,6'd53,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd68: Enemy_img = 4'd13;
//6'd47,6'd48,6'd51,6'd52,6'd53,6'd56,6'd59,6'd60,6'd61,6'd63,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd50,6'd54,6'd55,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd61,6'd69: Enemy_img = 4'd13;
//6'd46,6'd47,6'd52,6'd53,6'd54,6'd56,6'd59,6'd60,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd50,6'd51,6'd55,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd61,6'd69: Enemy_img = 4'd13;
//6'd46,6'd47,6'd49,6'd52,6'd53,6'd55,6'd59,6'd60,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd51,6'd54,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd60,6'd71: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd49,6'd52,6'd53,6'd55,6'd58,6'd59,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd43,6'd44,6'd51,6'd54,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd60,6'd71,6'd72: Enemy_img = 4'd13;
//6'd45,6'd46,6'd48,6'd53,6'd58,6'd59,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd77,6'd78: Enemy_img = 4'd14;
//6'd49,6'd51,6'd52,6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd72: Enemy_img = 4'd13;
//6'd48,6'd53,6'd54,6'd57,6'd58,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd49,6'd51,6'd52,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd13;
//6'd53,6'd57,6'd58,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd52,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd72: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd73: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd72: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd73: Enemy_img = 4'd14;
//6'd52,6'd53,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd71: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd52,6'd67,6'd68,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd71: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd52,6'd66,6'd67,6'd68,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd70: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd61,6'd62,6'd63,6'd68,6'd69,6'd71: Enemy_img = 4'd14;
//6'd65,6'd66,6'd67,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd70: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd61,6'd62,6'd68,6'd69,6'd71: Enemy_img = 4'd14;
//6'd67,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd70: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd71: Enemy_img = 4'd14;
//6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd56,6'd57,6'd60: Enemy_img = 4'd14;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd56,6'd57: Enemy_img = 4'd14;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55: Enemy_img = 4'd13;
//6'd52,6'd53,6'd56,6'd57: Enemy_img = 4'd14;
//6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd13;
//6'd52,6'd53,6'd55,6'd56: Enemy_img = 4'd14;
//6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd55,6'd56: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd51,6'd52,6'd54,6'd55: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd51,6'd52,6'd54,6'd55: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd54: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd48: Enemy_img = 4'd14;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd48: Enemy_img = 4'd14;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd14;
//6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd14;
//6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd59,6'd60,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd57,6'd58,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd74,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd70,6'd73,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd70,6'd73,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd72: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd48,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd66,6'd67,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd63,6'd71,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd72,6'd73: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd70,6'd71: Enemy_img = 4'd13;
//6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd74,6'd75: Enemy_img = 4'd14;
//6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd69,6'd70,6'd73: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd67,6'd68,6'd74: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd66,6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd67,6'd68,6'd69,6'd73,6'd74: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd72: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd52,6'd53,6'd57,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd71: Enemy_img = 4'd13;
//6'd52,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd73: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd68,6'd70,6'd74: Enemy_img = 4'd13;
//6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd69,6'd71,6'd72,6'd75,6'd76: Enemy_img = 4'd14;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd70,6'd71,6'd72,6'd75: Enemy_img = 4'd13;
//6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd73,6'd76,6'd77: Enemy_img = 4'd14;
//6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd70,6'd71,6'd74: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd67,6'd72,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd66: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65: Enemy_img = 4'd10;
//6'd68,6'd69,6'd70,6'd73: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd49,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd65,6'd66,6'd67: Enemy_img = 4'd9;
//6'd64: Enemy_img = 4'd10;
//6'd69: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd49,6'd55,6'd60,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd9;
//6'd71: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd49,6'd56,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd71: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd54,6'd55,6'd58,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd65,6'd66,6'd68,6'd71: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd54,6'd55,6'd58,6'd61,6'd62,6'd63,6'd64,6'd67,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd50,6'd53,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd71: Enemy_img = 4'd13;
//6'd51,6'd52,6'd54,6'd55,6'd58,6'd59,6'd60,6'd67,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84: Enemy_img = 4'd14;
//6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd66: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65: Enemy_img = 4'd10;
//6'd68,6'd71: Enemy_img = 4'd13;
//6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd54,6'd55,6'd58,6'd59,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd43,6'd50,6'd53,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd65,6'd66,6'd67: Enemy_img = 4'd9;
//6'd64: Enemy_img = 4'd10;
//6'd69,6'd72: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd57,6'd58,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd42,6'd50,6'd53,6'd54,6'd55,6'd60,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd9;
//6'd69: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd42,6'd50,6'd55,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd72: Enemy_img = 4'd13;
//6'd35,6'd37,6'd38,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd39,6'd40,6'd41,6'd50,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd65,6'd66,6'd68,6'd69,6'd72: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd40,6'd43,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd67,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd36,6'd39,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd70,6'd73: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd67,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd44,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd66: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65: Enemy_img = 4'd10;
//6'd68,6'd69,6'd73: Enemy_img = 4'd13;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd32,6'd33,6'd35,6'd42,6'd44,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd65,6'd66,6'd67: Enemy_img = 4'd9;
//6'd64: Enemy_img = 4'd10;
//6'd71,6'd74: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd69,6'd70,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd34,6'd35,6'd43,6'd45,6'd46,6'd47,6'd48,6'd53,6'd60,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd9;
//6'd69,6'd71,6'd72,6'd75: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd70,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd36,6'd37,6'd41,6'd42,6'd43,6'd48,6'd52,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd71,6'd72,6'd73,6'd76: Enemy_img = 4'd13;
//6'd40,6'd42,6'd43,6'd46,6'd47,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd70,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd41,6'd44,6'd48,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd65,6'd66,6'd67,6'd71,6'd72,6'd73,6'd77: Enemy_img = 4'd13;
//6'd42,6'd43,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd70,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd44,6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd76: Enemy_img = 4'd13;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd41,6'd42,6'd45,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd69,6'd74,6'd75: Enemy_img = 4'd13;
//6'd44,6'd47,6'd48,6'd49,6'd51,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd70,6'd71,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd42,6'd43,6'd45,6'd50,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd72,6'd73: Enemy_img = 4'd13;
//6'd45,6'd48,6'd49,6'd51,6'd52,6'd53,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd43,6'd44,6'd46,6'd50,6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd70,6'd71: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd50,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd49,6'd50,6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd70,6'd71: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd68,6'd69,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd46,6'd47,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd72: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd47,6'd48,6'd50,6'd51,6'd57,6'd58,6'd59,6'd60,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd74,6'd75: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd60,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd79: Enemy_img = 4'd14;
//6'd48,6'd55,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd76: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//6'd50,6'd55,6'd56,6'd57,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd48,6'd50,6'd51,6'd55,6'd60,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd54,6'd55,6'd56,6'd57,6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd78: Enemy_img = 4'd14;
//6'd48,6'd49,6'd52,6'd53,6'd58,6'd60,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd55,6'd56,6'd57,6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd53,6'd54,6'd58,6'd60,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd56,6'd57,6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd54,6'd55,6'd58,6'd60,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd57,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd55,6'd56,6'd58,6'd59,6'd60,6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd57,6'd58,6'd59,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd54,6'd56,6'd60,6'd73,6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd58,6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd54,6'd56,6'd57,6'd59,6'd73,6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd64,6'd77: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd58,6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69,6'd70,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd54,6'd55,6'd57,6'd59,6'd72,6'd73,6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd57,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd14;
//6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd14;
//6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66,6'd68: Enemy_img = 4'd14;
//6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66,6'd68: Enemy_img = 4'd14;
//6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd13;
//6'd47,6'd50,6'd51,6'd52,6'd59,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd13;
//6'd47,6'd50,6'd51,6'd53,6'd59,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd52,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd48,6'd51,6'd53,6'd57,6'd58,6'd59,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd52,6'd55,6'd58,6'd60,6'd61: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd48,6'd51,6'd53,6'd54,6'd56,6'd57,6'd59,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd53,6'd55,6'd57,6'd58: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd52,6'd54,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd52,6'd54,6'd57,6'd62,6'd63: Enemy_img = 4'd14;
//6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd54,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd53,6'd55,6'd56,6'd57,6'd58,6'd62,6'd63: Enemy_img = 4'd14;
//6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd59: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd62: Enemy_img = 4'd14;
//6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd54,6'd55,6'd57,6'd58,6'd59: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd56: Enemy_img = 4'd14;
//6'd35,6'd36: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd55,6'd57,6'd58,6'd61: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd54,6'd56,6'd59,6'd60,6'd62,6'd63: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd55,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd51,6'd54,6'd56,6'd57,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd33,6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd51,6'd55,6'd56,6'd57,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd33: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd32: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66: Enemy_img = 4'd13;
//6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd59,6'd61,6'd62,6'd63: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd65: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd61,6'd62: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd60,6'd61,6'd62: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59: Enemy_img = 4'd9;
//6'd61,6'd64: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60: Enemy_img = 4'd9;
//6'd56,6'd57: Enemy_img = 4'd10;
//6'd64: Enemy_img = 4'd13;
//6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56: Enemy_img = 4'd9;
//6'd57: Enemy_img = 4'd10;
//6'd65: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55: Enemy_img = 4'd9;
//6'd58,6'd59,6'd60,6'd62,6'd65: Enemy_img = 4'd13;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd61,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd45,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd66,6'd67: Enemy_img = 4'd13;
//6'd43,6'd44,6'd49,6'd50,6'd51,6'd52,6'd61,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd63: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd56,6'd57,6'd58,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd9;
//6'd59,6'd60: Enemy_img = 4'd10;
//6'd54,6'd64,6'd67: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd55,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd61,6'd62: Enemy_img = 4'd9;
//6'd59,6'd60: Enemy_img = 4'd10;
//6'd64,6'd65,6'd68: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd43,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58: Enemy_img = 4'd9;
//6'd64,6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd13;
//6'd42,6'd45,6'd49,6'd50,6'd53,6'd54,6'd67,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd43,6'd44,6'd46,6'd47,6'd48,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd70,6'd71: Enemy_img = 4'd13;
//6'd42,6'd43,6'd47,6'd49,6'd50,6'd53,6'd54,6'd63,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd48,6'd51,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd61,6'd65,6'd68,6'd73,6'd74: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd50,6'd53,6'd54,6'd60,6'd66,6'd67,6'd69,6'd70,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd45,6'd49,6'd51,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd9;
//6'd62: Enemy_img = 4'd10;
//6'd57,6'd68,6'd69,6'd70,6'd75: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd47,6'd48,6'd53,6'd54,6'd58,6'd59,6'd66,6'd67,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd49,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64: Enemy_img = 4'd9;
//6'd60,6'd61,6'd62: Enemy_img = 4'd10;
//6'd56,6'd67,6'd69,6'd70,6'd71,6'd74: Enemy_img = 4'd13;
//6'd45,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd57,6'd68,6'd72,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd46,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60: Enemy_img = 4'd9;
//6'd61,6'd62: Enemy_img = 4'd10;
//6'd69,6'd70,6'd73,6'd74: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd67,6'd68,6'd71,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd41,6'd47,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd68,6'd69,6'd72,6'd73: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd66,6'd67,6'd70,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd14;
//6'd39,6'd47,6'd52,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd72: Enemy_img = 4'd13;
//6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd67,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd14;
//6'd39,6'd47,6'd52,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd64,6'd65,6'd66,6'd71: Enemy_img = 4'd13;
//6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd39,6'd45,6'd46,6'd47,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd64,6'd65,6'd66,6'd70: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd41,6'd42,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd39,6'd43,6'd44,6'd45: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd71,6'd72: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd69: Enemy_img = 4'd14;
//6'd38,6'd39,6'd42,6'd43,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd68,6'd73,6'd75,6'd76,6'd77: Enemy_img = 4'd13;
//6'd35,6'd36,6'd38,6'd44,6'd45,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd69,6'd70,6'd71,6'd72,6'd74,6'd78: Enemy_img = 4'd14;
//6'd37,6'd39,6'd40,6'd42,6'd43,6'd46,6'd47,6'd51,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd46,6'd48,6'd49,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd14;
//6'd34,6'd37,6'd41,6'd44,6'd45,6'd47,6'd50,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd42,6'd48,6'd49,6'd50,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd79: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd46,6'd47,6'd48,6'd49,6'd52,6'd60,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd14;
//6'd34,6'd35,6'd41,6'd42,6'd43,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd80: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd64,6'd65,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd81: Enemy_img = 4'd14;
//6'd34,6'd35,6'd41,6'd44,6'd45,6'd51,6'd57,6'd62,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd80: Enemy_img = 4'd13;
//6'd30,6'd40,6'd43,6'd44,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd62,6'd64,6'd65,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd81: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd45,6'd46,6'd51,6'd56,6'd60,6'd61,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd81: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd49,6'd50,6'd52,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd64,6'd65,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd82: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd51,6'd55,6'd59,6'd60,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd81: Enemy_img = 4'd13;
//6'd52,6'd53,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd65,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd82: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd54,6'd59,6'd63,6'd77,6'd78,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd81,6'd82: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd79,6'd80: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd58,6'd59,6'd63,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd59,6'd62,6'd66,6'd67,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd80: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd58,6'd60,6'd61,6'd63,6'd64,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd60,6'd61,6'd63,6'd66,6'd67,6'd69,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd50,6'd51,6'd53,6'd54,6'd58,6'd59,6'd62,6'd64,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd13;
//6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd67,6'd68,6'd70,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd57,6'd62,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd13;
//6'd59,6'd60,6'd61,6'd62,6'd67,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd52,6'd56,6'd57,6'd58,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70: Enemy_img = 4'd13;
//6'd54,6'd55,6'd62,6'd63,6'd64,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//6'd52,6'd53,6'd58,6'd59,6'd60,6'd61,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd70: Enemy_img = 4'd13;
//6'd55,6'd56,6'd63,6'd64,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd61,6'd62,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd70: Enemy_img = 4'd13;
//6'd55,6'd56,6'd58,6'd59,6'd64,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd75: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd60,6'd62,6'd63,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd71: Enemy_img = 4'd13;
//6'd56,6'd57,6'd59,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd75: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd71: Enemy_img = 4'd13;
//6'd56,6'd57,6'd59,6'd68,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd60,6'd61,6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd13;
//6'd69,6'd70,6'd71,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd70,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd70,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd13;
//6'd71,6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd13;
//6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd72,6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd13;
//6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd13;
//6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd74,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd75,6'd76,6'd78,6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd13;
//6'd76,6'd77: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd13;
//6'd77: Enemy_img = 4'd14;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd13;
//6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd13;
//6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd13;
//6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd48: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd45,6'd46,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd47: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd41,6'd42,6'd45,6'd46: Enemy_img = 4'd13;
//6'd37,6'd40,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd39,6'd40,6'd42,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd13;
//6'd34,6'd38,6'd41,6'd43,6'd44,6'd49,6'd50,6'd81: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd40,6'd41,6'd43,6'd47,6'd48: Enemy_img = 4'd13;
//6'd35,6'd39,6'd42,6'd44,6'd45,6'd46,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd30,6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd41,6'd42,6'd48,6'd50: Enemy_img = 4'd13;
//6'd32,6'd33,6'd36,6'd40,6'd43,6'd44,6'd45,6'd46,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd31: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd42,6'd47,6'd48,6'd50: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd37,6'd41,6'd44,6'd49,6'd51,6'd52,6'd53,6'd54,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd45,6'd52,6'd53,6'd54,6'd55,6'd56,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd30: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd45,6'd46,6'd49,6'd55,6'd57: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd44,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd51,6'd52,6'd57: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd29: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd48,6'd49,6'd50,6'd57: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd46,6'd47,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd53,6'd54,6'd55,6'd57: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd43,6'd50,6'd51,6'd52,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd28: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd51,6'd53,6'd54,6'd55: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd44,6'd48,6'd49,6'd50,6'd52,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd51,6'd53,6'd54,6'd55: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd47,6'd49,6'd50,6'd52,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd53,6'd54,6'd55,6'd57: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd52,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd26,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd54,6'd55,6'd58: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd26,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53: Enemy_img = 4'd9;
//6'd50,6'd59: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54: Enemy_img = 4'd9;
//6'd51: Enemy_img = 4'd10;
//6'd60,6'd61: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd57,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd25,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52: Enemy_img = 4'd10;
//6'd57: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd56,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd25,6'd31,6'd32,6'd33,6'd34,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51: Enemy_img = 4'd9;
//6'd53,6'd54,6'd55,6'd58,6'd59,6'd63,6'd64,6'd65: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd60,6'd61,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd57: Enemy_img = 4'd9;
//6'd52,6'd53,6'd54,6'd60,6'd66,6'd71: Enemy_img = 4'd13;
//6'd25,6'd37,6'd38,6'd39,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd61,6'd62,6'd63,6'd72,6'd73,6'd74,6'd77,6'd78: Enemy_img = 4'd14;
//6'd24,6'd26,6'd27,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58: Enemy_img = 4'd9;
//6'd55: Enemy_img = 4'd10;
//6'd51,6'd52,6'd60,6'd61,6'd62,6'd63,6'd71: Enemy_img = 4'd13;
//6'd38,6'd43,6'd44,6'd45,6'd46,6'd47,6'd53,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd24,6'd39,6'd40,6'd41,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56: Enemy_img = 4'd10;
//6'd51,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd71: Enemy_img = 4'd13;
//6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd60,6'd63,6'd64,6'd69,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd38,6'd39,6'd41,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55: Enemy_img = 4'd9;
//6'd51,6'd58,6'd59,6'd62,6'd66,6'd67,6'd68: Enemy_img = 4'd13;
//6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd60,6'd61,6'd63,6'd64,6'd65,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54: Enemy_img = 4'd9;
//6'd50,6'd57,6'd58,6'd64,6'd67,6'd70: Enemy_img = 4'd13;
//6'd39,6'd40,6'd49,6'd51,6'd65,6'd66,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62: Enemy_img = 4'd9;
//6'd56,6'd67,6'd70: Enemy_img = 4'd13;
//6'd40,6'd42,6'd43,6'd44,6'd45,6'd50,6'd51,6'd57,6'd58,6'd65,6'd66,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd41,6'd46,6'd47,6'd53,6'd54,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd9;
//6'd59,6'd60: Enemy_img = 4'd10;
//6'd55,6'd66,6'd67,6'd70: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd56,6'd57,6'd64,6'd65,6'd68,6'd71,6'd72,6'd73,6'd77,6'd78: Enemy_img = 4'd14;
//6'd48,6'd53,6'd54,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd9;
//6'd59,6'd60: Enemy_img = 4'd10;
//6'd55,6'd62,6'd63,6'd64,6'd67,6'd69,6'd75,6'd76: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd52,6'd56,6'd65,6'd66,6'd77,6'd78,6'd80: Enemy_img = 4'd14;
//6'd49,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59: Enemy_img = 4'd9;
//6'd54,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd71,6'd72: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd47,6'd48,6'd51,6'd52,6'd53,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd49,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd80: Enemy_img = 4'd13;
//6'd45,6'd46,6'd48,6'd52,6'd53,6'd54,6'd55,6'd56,6'd62,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd47,6'd49,6'd50,6'd58,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd64,6'd65,6'd68,6'd81: Enemy_img = 4'd13;
//6'd41,6'd45,6'd46,6'd47,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd82,6'd83: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd51,6'd58,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd65,6'd82,6'd83: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd84: Enemy_img = 4'd14;
//6'd44,6'd45,6'd51,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd83,6'd84: Enemy_img = 4'd13;
//6'd41,6'd42,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd41,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd42,6'd43,6'd47,6'd52,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82: Enemy_img = 4'd14;
//6'd41,6'd42,6'd47,6'd48,6'd52,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd67,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd47,6'd48,6'd52,6'd65,6'd66,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd62,6'd63,6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd40,6'd46,6'd47,6'd52,6'd60,6'd64,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd62,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd40,6'd45,6'd46,6'd52,6'd58,6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd13;
//6'd39,6'd40,6'd43,6'd46,6'd47,6'd50,6'd51,6'd58,6'd61,6'd62,6'd64,6'd65,6'd68,6'd69,6'd70,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd41,6'd44,6'd45,6'd48,6'd49,6'd52,6'd55,6'd56,6'd57,6'd59,6'd63,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd39,6'd40,6'd43,6'd46,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd64,6'd65,6'd69,6'd70,6'd71,6'd73,6'd74,6'd78,6'd79: Enemy_img = 4'd14;
//6'd41,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd59,6'd62,6'd63,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd39,6'd40,6'd48,6'd49,6'd50,6'd52,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd79,6'd80: Enemy_img = 4'd14;
//6'd41,6'd45,6'd46,6'd47,6'd51,6'd53,6'd54,6'd59,6'd63,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd13;
//6'd38,6'd39,6'd42,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd60,6'd61,6'd64,6'd67,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd40,6'd41,6'd43,6'd44,6'd54,6'd55,6'd58,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54,6'd57,6'd60,6'd61,6'd62,6'd68,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd40,6'd41,6'd46,6'd47,6'd55,6'd56,6'd58,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd47,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd41,6'd45,6'd46,6'd48,6'd49,6'd50,6'd55,6'd58,6'd63,6'd68,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd45,6'd46,6'd52,6'd53,6'd62,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd13;
//6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd68,6'd69,6'd70,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd38,6'd39,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd13;
//6'd37,6'd38,6'd40,6'd41,6'd42,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd39,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd52,6'd53,6'd56,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd80: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd61,6'd62,6'd65,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd58,6'd59,6'd60,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd81: Enemy_img = 4'd13;
//6'd36,6'd62,6'd63,6'd66,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd59,6'd60,6'd61,6'd67,6'd68,6'd73,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd82: Enemy_img = 4'd13;
//6'd35,6'd63,6'd64,6'd67,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd83: Enemy_img = 4'd13;
//6'd63,6'd64,6'd65,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd13;
//6'd64,6'd65,6'd81,6'd82,6'd83,6'd85,6'd86: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd63,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85: Enemy_img = 4'd13;
//6'd82,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd14;
//6'd61,6'd62,6'd63,6'd64,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86: Enemy_img = 4'd13;
//6'd83,6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd62,6'd63,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87: Enemy_img = 4'd13;
//6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd14;
//6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88: Enemy_img = 4'd13;
//6'd85,6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89: Enemy_img = 4'd13;
//6'd86,6'd87,6'd88,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90: Enemy_img = 4'd13;
//6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91: Enemy_img = 4'd13;
//6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92: Enemy_img = 4'd13;
//6'd91: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93: Enemy_img = 4'd13;
//6'd92: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd38,6'd39,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd13;
//6'd34,6'd35,6'd38,6'd39,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd13;
//6'd33,6'd34,6'd38,6'd39,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd38,6'd39,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd38,6'd39,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd40,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd36,6'd37: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd34,6'd35,6'd38,6'd39,6'd40,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd39: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd39: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd37,6'd40,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd34,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd39,6'd41,6'd42: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd34,6'd35,6'd39,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49: Enemy_img = 4'd13;
//6'd27,6'd28,6'd31,6'd32,6'd33,6'd36,6'd40,6'd44,6'd45,6'd46,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd13;
//6'd29,6'd30,6'd34,6'd35,6'd36,6'd44,6'd45,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28,6'd34,6'd39,6'd40,6'd41,6'd44,6'd45,6'd48,6'd50: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd37,6'd38,6'd42,6'd43,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd43,6'd44,6'd47,6'd48: Enemy_img = 4'd13;
//6'd26,6'd27,6'd33,6'd39,6'd40,6'd41,6'd42,6'd46,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd36,6'd42,6'd46,6'd47,6'd48,6'd49,6'd51,6'd66: Enemy_img = 4'd13;
//6'd29,6'd30,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd14;
//6'd25: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd41,6'd45,6'd48,6'd49,6'd52,6'd53,6'd64,6'd65: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd39,6'd40,6'd44,6'd46,6'd47,6'd50,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd43,6'd45,6'd48,6'd49,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd67: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd42,6'd44,6'd46,6'd47,6'd50,6'd57,6'd58,6'd59,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74: Enemy_img = 4'd14;
//6'd23,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd43,6'd45,6'd46,6'd67: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd36,6'd37,6'd42,6'd44,6'd47,6'd51,6'd52,6'd53,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd23,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50: Enemy_img = 4'd9;
//6'd45,6'd46,6'd52,6'd63,6'd64,6'd67: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd23,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49: Enemy_img = 4'd9;
//6'd47: Enemy_img = 4'd10;
//6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd67,6'd73,6'd74,6'd77,6'd78: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd60,6'd65,6'd68,6'd69,6'd70,6'd71,6'd75,6'd79,6'd80: Enemy_img = 4'd14;
//6'd23,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd54,6'd55: Enemy_img = 4'd9;
//6'd47: Enemy_img = 4'd10;
//6'd50,6'd51,6'd57,6'd58,6'd59,6'd63,6'd64,6'd65,6'd67,6'd72,6'd73,6'd79,6'd80: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd60,6'd61,6'd62,6'd68,6'd69,6'd71,6'd74,6'd75,6'd76,6'd78,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55: Enemy_img = 4'd9;
//6'd46,6'd47: Enemy_img = 4'd10;
//6'd50,6'd51,6'd58,6'd59,6'd62,6'd64,6'd65,6'd67,6'd68,6'd81,6'd82,6'd83: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd57,6'd61,6'd63,6'd66,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd23: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd54: Enemy_img = 4'd9;
//6'd52,6'd53: Enemy_img = 4'd10;
//6'd49,6'd56,6'd57,6'd64,6'd65,6'd67,6'd70,6'd71: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd50,6'd63,6'd66,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd23,6'd39: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd59,6'd60,6'd61: Enemy_img = 4'd9;
//6'd52,6'd53: Enemy_img = 4'd10;
//6'd49,6'd55,6'd56,6'd69: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd50,6'd63,6'd64,6'd65,6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd81,6'd82: Enemy_img = 4'd14;
//6'd23,6'd39,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd59: Enemy_img = 4'd9;
//6'd58: Enemy_img = 4'd10;
//6'd55,6'd62,6'd63,6'd64: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd49,6'd56,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd23,6'd39,6'd46,6'd47,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd9;
//6'd58,6'd59: Enemy_img = 4'd10;
//6'd49,6'd54,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd55,6'd56,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd23,6'd39,6'd47,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd9;
//6'd49,6'd54,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd50,6'd55,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd23,6'd39,6'd52,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd9;
//6'd54,6'd60,6'd65: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd55,6'd61,6'd62,6'd63,6'd64,6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd23,6'd32,6'd38,6'd39,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd9;
//6'd54,6'd60,6'd68: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd36,6'd41,6'd42,6'd43,6'd49,6'd50,6'd51,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd23,6'd29,6'd30,6'd37,6'd38,6'd39,6'd46,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd68,6'd69: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd38,6'd39,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd23,6'd28,6'd37,6'd40,6'd44,6'd47,6'd48,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd70,6'd71: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd23,6'd27,6'd40,6'd41,6'd42,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd72,6'd73,6'd74: Enemy_img = 4'd13;
//6'd24,6'd25,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd23,6'd26,6'd50,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd13;
//6'd24,6'd40,6'd41,6'd42,6'd43,6'd44,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd23,6'd25,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd67,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd23,6'd24,6'd45,6'd49,6'd53,6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80,6'd81: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd64,6'd65,6'd67,6'd68,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd23,6'd41,6'd42,6'd43,6'd44,6'd45,6'd54,6'd62,6'd66,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83: Enemy_img = 4'd13;
//6'd42,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd64,6'd67,6'd68,6'd69,6'd70,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd43,6'd44,6'd46,6'd47,6'd62,6'd65,6'd66,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85,6'd86: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd62,6'd64,6'd65,6'd68,6'd71,6'd72,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49,6'd50,6'd55,6'd60,6'd61,6'd66,6'd67,6'd69,6'd70,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88: Enemy_img = 4'd13;
//6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd57,6'd61,6'd64,6'd65,6'd68,6'd70,6'd74,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd45,6'd50,6'd55,6'd59,6'd60,6'd62,6'd66,6'd67,6'd69,6'd71,6'd72,6'd73,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89,6'd90: Enemy_img = 4'd13;
//6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd62,6'd64,6'd65,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd45,6'd50,6'd58,6'd59,6'd66,6'd67,6'd68,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92,6'd93: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd94,6'd95: Enemy_img = 4'd14;
//6'd50,6'd56,6'd57,6'd67,6'd68,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd69,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd49,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd96,6'd97: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd62,6'd64,6'd65,6'd66,6'd91,6'd92,6'd93,6'd94,6'd95,6'd98: Enemy_img = 4'd14;
//6'd44,6'd49,6'd52,6'd55,6'd60,6'd61,6'd63,6'd67,6'd68,6'd69,6'd70,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd99,6'd100: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd71,6'd72,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd44,6'd45,6'd49,6'd51,6'd52,6'd60,6'd65,6'd66,6'd67,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72,6'd101,6'd102: Enemy_img = 4'd13;
//6'd44,6'd48,6'd68,6'd69,6'd73,6'd74,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd45,6'd46,6'd50,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd44,6'd45,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd101,6'd102: Enemy_img = 4'd14;
//6'd46,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd51,6'd52,6'd58,6'd59,6'd60,6'd61,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd72,6'd73: Enemy_img = 4'd14;
//6'd46,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd47,6'd52,6'd53,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd48,6'd49: Enemy_img = 4'd14;
//6'd46,6'd47,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd14;
//6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd14;
//6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92: Enemy_img = 4'd13;
//6'd93: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91: Enemy_img = 4'd13;
//6'd92: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90: Enemy_img = 4'd13;
//6'd91: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89: Enemy_img = 4'd13;
//6'd87,6'd88,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88: Enemy_img = 4'd13;
//6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87: Enemy_img = 4'd13;
//6'd85,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86: Enemy_img = 4'd13;
//6'd84,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85: Enemy_img = 4'd13;
//6'd82,6'd83,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd13;
//6'd81,6'd82,6'd83,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd61,6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd83: Enemy_img = 4'd13;
//6'd63,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd82: Enemy_img = 4'd13;
//6'd62,6'd65,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd81: Enemy_img = 4'd13;
//6'd61,6'd62,6'd64,6'd65,6'd66,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd59,6'd60,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd80: Enemy_img = 4'd13;
//6'd34,6'd35,6'd60,6'd61,6'd63,6'd64,6'd65,6'd74,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd59,6'd66,6'd67,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd79: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd59,6'd60,6'd62,6'd63,6'd64,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd58,6'd65,6'd66,6'd67,6'd68,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd58,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd75: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd74: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd71: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd60,6'd70: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd69: Enemy_img = 4'd13;
//6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72,6'd76,6'd77: Enemy_img = 4'd14;
//6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd68: Enemy_img = 4'd13;
//6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd76,6'd77: Enemy_img = 4'd14;
//6'd73,6'd74,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd62,6'd65,6'd66,6'd67: Enemy_img = 4'd13;
//6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd56,6'd57,6'd58,6'd68,6'd69,6'd70,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd72,6'd73,6'd75,6'd78,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd66: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd60,6'd61,6'd67,6'd68,6'd69,6'd73,6'd75,6'd76,6'd81: Enemy_img = 4'd14;
//6'd71,6'd72,6'd74,6'd77,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd54,6'd55,6'd58,6'd61,6'd81,6'd82: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd68,6'd72,6'd75,6'd76,6'd80: Enemy_img = 4'd14;
//6'd67,6'd70,6'd71,6'd73,6'd74,6'd77,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd54,6'd60,6'd61,6'd62,6'd63,6'd80,6'd81: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd79,6'd82,6'd83: Enemy_img = 4'd14;
//6'd67,6'd73,6'd74,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd56,6'd59,6'd60,6'd61,6'd62,6'd79,6'd80: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd58,6'd63,6'd64,6'd65,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd68,6'd69,6'd74,6'd77,6'd78,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd9;
//6'd51,6'd53,6'd54,6'd59,6'd60,6'd61,6'd79: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd55,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd80,6'd81: Enemy_img = 4'd14;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd9;
//6'd53,6'd54,6'd55,6'd59,6'd60: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd72,6'd75,6'd79,6'd80: Enemy_img = 4'd14;
//6'd71,6'd73,6'd74,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd9;
//6'd49,6'd53,6'd54,6'd60,6'd61: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd52,6'd55,6'd62,6'd63,6'd64,6'd65,6'd66,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd79: Enemy_img = 4'd14;
//6'd73,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd9;
//6'd58,6'd59: Enemy_img = 4'd10;
//6'd49,6'd52,6'd53,6'd61,6'd62: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd54,6'd55,6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd68,6'd69,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60: Enemy_img = 4'd9;
//6'd58,6'd59: Enemy_img = 4'd10;
//6'd48,6'd51,6'd55,6'd63,6'd64: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd65,6'd66,6'd67,6'd75,6'd76: Enemy_img = 4'd14;
//6'd69,6'd70,6'd71,6'd72,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd59,6'd60: Enemy_img = 4'd9;
//6'd47,6'd51,6'd55,6'd56: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd50,6'd57,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd61,6'd62,6'd69,6'd73,6'd74,6'd75,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd60: Enemy_img = 4'd9;
//6'd40,6'd41,6'd42,6'd43,6'd46,6'd50,6'd56: Enemy_img = 4'd13;
//6'd39,6'd44,6'd45,6'd49,6'd57,6'd58,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd9;
//6'd54: Enemy_img = 4'd10;
//6'd57: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd42,6'd47,6'd48,6'd50,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd75: Enemy_img = 4'd14;
//6'd70,6'd74,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55: Enemy_img = 4'd9;
//6'd53,6'd54: Enemy_img = 4'd10;
//6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd58,6'd59,6'd60: Enemy_img = 4'd13;
//6'd38,6'd39,6'd42,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72: Enemy_img = 4'd14;
//6'd70,6'd73,6'd74,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd55,6'd56: Enemy_img = 4'd9;
//6'd54: Enemy_img = 4'd10;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd60: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd42,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd74: Enemy_img = 4'd14;
//6'd57,6'd58,6'd72,6'd73,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd55,6'd56: Enemy_img = 4'd9;
//6'd43,6'd44,6'd45,6'd46,6'd51,6'd52: Enemy_img = 4'd13;
//6'd23,6'd24,6'd37,6'd38,6'd39,6'd40,6'd42,6'd53,6'd60,6'd61,6'd62,6'd63,6'd73,6'd74: Enemy_img = 4'd14;
//6'd57,6'd58,6'd71,6'd72,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49: Enemy_img = 4'd9;
//6'd50: Enemy_img = 4'd10;
//6'd41,6'd52,6'd53: Enemy_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd37,6'd38,6'd39,6'd40,6'd43,6'd44,6'd45,6'd46,6'd54,6'd59,6'd60,6'd61,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd9;
//6'd49,6'd50: Enemy_img = 4'd10;
//6'd38,6'd39,6'd41,6'd44,6'd45,6'd46,6'd53,6'd54,6'd55: Enemy_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd37,6'd40,6'd43,6'd56,6'd57,6'd58,6'd59,6'd60,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd76: Enemy_img = 4'd14;
//6'd62,6'd63,6'd71,6'd72,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd9;
//6'd50: Enemy_img = 4'd10;
//6'd26,6'd36,6'd37,6'd38,6'd39,6'd42,6'd46,6'd47,6'd48,6'd56: Enemy_img = 4'd13;
//6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd43,6'd44,6'd45,6'd57,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd76: Enemy_img = 4'd14;
//6'd61,6'd62,6'd71,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd9;
//6'd27,6'd28,6'd29,6'd38,6'd39,6'd40,6'd42: Enemy_img = 4'd13;
//6'd25,6'd26,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd56,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd76: Enemy_img = 4'd14;
//6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd70,6'd71,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd45: Enemy_img = 4'd13;
//6'd25,6'd26,6'd32,6'd33,6'd40,6'd41,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd55,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd68,6'd69,6'd72,6'd73,6'd76: Enemy_img = 4'd14;
//6'd58,6'd62,6'd66,6'd67,6'd70,6'd71,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd38,6'd39: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd33,6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd75,6'd76: Enemy_img = 4'd14;
//6'd57,6'd61,6'd65,6'd66,6'd67,6'd68,6'd72,6'd74,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd33,6'd34,6'd38,6'd40: Enemy_img = 4'd13;
//6'd26,6'd27,6'd31,6'd32,6'd35,6'd36,6'd39,6'd41,6'd42,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd70,6'd71: Enemy_img = 4'd14;
//6'd57,6'd60,6'd64,6'd68,6'd69,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd33,6'd34,6'd39,6'd40,6'd44: Enemy_img = 4'd13;
//6'd26,6'd27,6'd30,6'd31,6'd32,6'd35,6'd36,6'd38,6'd41,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd74,6'd77: Enemy_img = 4'd14;
//6'd60,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd39,6'd43: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd44,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd65,6'd66,6'd67,6'd68,6'd69,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd70,6'd71,6'd73,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd35,6'd39,6'd42: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd33,6'd34,6'd36,6'd43,6'd46,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd47,6'd48,6'd61,6'd62,6'd64,6'd65,6'd73,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd41: Enemy_img = 4'd13;
//6'd28,6'd29,6'd35,6'd42,6'd45,6'd46,6'd47,6'd48,6'd55,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd61,6'd62,6'd65,6'd66,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd40: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd34,6'd37,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61,6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd34,6'd35,6'd39: Enemy_img = 4'd13;
//6'd29,6'd30,6'd33,6'd36,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd70,6'd71,6'd72,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd53,6'd68,6'd69,6'd73,6'd74,6'd76,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd38: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd35,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd53,6'd54,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd37: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd34,6'd38,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd73,6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd54,6'd76,6'd77,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd49,6'd50,6'd51,6'd52,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd79,6'd80: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd13;
//6'd30,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd81: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd35,6'd36,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd35,6'd37,6'd38,6'd39,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd40,6'd41,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd42,6'd43,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd46,6'd47,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd14;
//6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd13;
//6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd13;
//6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd13;
//6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd13;
//6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd13;
//6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd13;
//6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd13;
//6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd13;
//6'd71,6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd13;
//6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd70,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72: Enemy_img = 4'd13;
//6'd69,6'd70,6'd73,6'd74: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd13;
//6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd13;
//6'd66,6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd70: Enemy_img = 4'd13;
//6'd55,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd70: Enemy_img = 4'd13;
//6'd55,6'd57,6'd58,6'd64,6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd53,6'd54,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd69: Enemy_img = 4'd13;
//6'd55,6'd57,6'd58,6'd63,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd59,6'd60,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd69: Enemy_img = 4'd13;
//6'd54,6'd56,6'd57,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd52,6'd53,6'd58,6'd59,6'd60,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd69: Enemy_img = 4'd13;
//6'd54,6'd56,6'd57,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd52,6'd53,6'd58,6'd59,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd68: Enemy_img = 4'd13;
//6'd53,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd52,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd68: Enemy_img = 4'd13;
//6'd53,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd52,6'd73,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd51,6'd73,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd68,6'd69,6'd73: Enemy_img = 4'd14;
//6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd66,6'd67: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd68,6'd69,6'd72,6'd73,6'd78: Enemy_img = 4'd14;
//6'd71,6'd74,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd66,6'd79: Enemy_img = 4'd13;
//6'd48,6'd49,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd67,6'd68,6'd73,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd70,6'd71,6'd72,6'd74,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd66,6'd78: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd67,6'd68,6'd71,6'd73,6'd74,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd70,6'd72,6'd75,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd65,6'd78: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd66,6'd67,6'd71,6'd73,6'd74,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd69,6'd70,6'd72,6'd75,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd65,6'd78: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd66,6'd67,6'd70,6'd72,6'd73,6'd74,6'd79,6'd80: Enemy_img = 4'd14;
//6'd69,6'd71,6'd75,6'd76,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd64: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd63,6'd65,6'd66,6'd67,6'd70,6'd73,6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd69,6'd71,6'd72,6'd76,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd78,6'd79: Enemy_img = 4'd14;
//6'd68,6'd73,6'd74,6'd75,6'd76,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd63,6'd64,6'd68,6'd69,6'd70,6'd79: Enemy_img = 4'd14;
//6'd66,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd63,6'd64,6'd65,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd70,6'd77,6'd78,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd56,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd73,6'd74,6'd75,6'd76,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd54,6'd56,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd55,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd69,6'd70,6'd72,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd9;
//6'd51,6'd54,6'd60,6'd61: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd55,6'd56,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//6'd71,6'd76,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd9;
//6'd51,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd13;
//6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd71,6'd72,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59: Enemy_img = 4'd9;
//6'd60: Enemy_img = 4'd10;
//6'd54,6'd55,6'd56,6'd66: Enemy_img = 4'd13;
//6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd67,6'd68,6'd69,6'd70,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd72,6'd73,6'd75,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd9;
//6'd59,6'd60: Enemy_img = 4'd10;
//6'd54,6'd55,6'd56: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd63,6'd64,6'd73,6'd75,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63: Enemy_img = 4'd9;
//6'd54,6'd55,6'd57: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd56,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd76,6'd77,6'd80: Enemy_img = 4'd14;
//6'd74,6'd75,6'd79,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd54,6'd57,6'd58: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd59,6'd60,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd76,6'd77,6'd80: Enemy_img = 4'd14;
//6'd74,6'd75,6'd79,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56: Enemy_img = 4'd9;
//6'd51,6'd58,6'd59: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd73,6'd74,6'd77,6'd80: Enemy_img = 4'd14;
//6'd71,6'd72,6'd75,6'd76,6'd79,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd9;
//6'd51,6'd54,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd14;
//6'd69,6'd75,6'd79,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd59: Enemy_img = 4'd9;
//6'd57,6'd58: Enemy_img = 4'd10;
//6'd50,6'd54: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd14;
//6'd68,6'd75,6'd79,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60: Enemy_img = 4'd9;
//6'd57,6'd58: Enemy_img = 4'd10;
//6'd50,6'd53: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd54,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd61,6'd62,6'd67,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60: Enemy_img = 4'd9;
//6'd49,6'd55,6'd56: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd54,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd82,6'd83: Enemy_img = 4'd14;
//6'd67,6'd77,6'd79,6'd80,6'd81,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd9;
//6'd47,6'd55,6'd56: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd50,6'd51,6'd57,6'd58,6'd61,6'd62,6'd63,6'd68,6'd69,6'd70,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd66,6'd67,6'd71,6'd72,6'd73,6'd74,6'd78,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54: Enemy_img = 4'd9;
//6'd45,6'd49,6'd50,6'd51,6'd57,6'd58,6'd60,6'd61: Enemy_img = 4'd13;
//6'd43,6'd44,6'd48,6'd59,6'd62,6'd63,6'd66,6'd69,6'd70,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd65,6'd67,6'd68,6'd71,6'd75,6'd76,6'd77,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55: Enemy_img = 4'd9;
//6'd45,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd43,6'd44,6'd46,6'd62,6'd65,6'd66,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd64,6'd67,6'd71,6'd80,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd9;
//6'd54,6'd55,6'd56: Enemy_img = 4'd10;
//6'd45,6'd48,6'd49: Enemy_img = 4'd13;
//6'd43,6'd44,6'd47,6'd50,6'd51,6'd52,6'd62,6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd81,6'd87: Enemy_img = 4'd14;
//6'd59,6'd60,6'd64,6'd67,6'd70,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd9;
//6'd56: Enemy_img = 4'd10;
//6'd49,6'd52,6'd53: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd48,6'd50,6'd51,6'd61,6'd62,6'd64,6'd65,6'd66,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd82,6'd83,6'd87: Enemy_img = 4'd14;
//6'd59,6'd63,6'd67,6'd70,6'd71,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd49,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd70,6'd71,6'd74,6'd75,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd72,6'd73,6'd77,6'd78,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd64,6'd69,6'd70,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd48,6'd51,6'd52: Enemy_img = 4'd13;
//6'd43,6'd44,6'd47,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd49: Enemy_img = 4'd13;
//6'd43,6'd47,6'd48,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd70,6'd71: Enemy_img = 4'd14;
//6'd65,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd50: Enemy_img = 4'd13;
//6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd65,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd45,6'd48,6'd49,6'd50,6'd55,6'd56,6'd66,6'd67: Enemy_img = 4'd14;
//6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd48,6'd49,6'd50,6'd53,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd46,6'd48,6'd52: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd47,6'd49,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65: Enemy_img = 4'd14;
//6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd43,6'd46,6'd48,6'd51: Enemy_img = 4'd13;
//6'd32,6'd33,6'd41,6'd42,6'd44,6'd47,6'd49,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd48,6'd49,6'd51: Enemy_img = 4'd13;
//6'd33,6'd34,6'd41,6'd44,6'd45,6'd46,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd45,6'd50: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd40,6'd41,6'd44,6'd46,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd45,6'd47,6'd50: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd49,6'd50: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd45,6'd47,6'd48,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd49: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd45,6'd47,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd46,6'd49: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd44,6'd45,6'd47,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd45,6'd48: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd44,6'd46,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd48: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd43,6'd44,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd49,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd63: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd58,6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd58,6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62,6'd74: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd68,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd47,6'd52,6'd53,6'd54,6'd67,6'd69,6'd71,6'd72,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62,6'd74: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd68,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd47,6'd52,6'd53,6'd67,6'd69,6'd70,6'd72,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62,6'd74: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67,6'd68,6'd69,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd47,6'd52,6'd53,6'd66,6'd70,6'd72,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62,6'd74: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd69,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd47,6'd52,6'd66,6'd67,6'd68,6'd70,6'd71,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62,6'd74: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67,6'd69,6'd70,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd47,6'd66,6'd68,6'd71,6'd72,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62: Enemy_img = 4'd13;
//6'd48,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67,6'd69,6'd70,6'd71,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd47,6'd66,6'd68,6'd72,6'd73,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd62: Enemy_img = 4'd13;
//6'd48,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67,6'd69,6'd70,6'd71,6'd72,6'd76: Enemy_img = 4'd14;
//6'd47,6'd66,6'd68,6'd73,6'd74,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67: Enemy_img = 4'd14;
//6'd47,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd47,6'd66,6'd71,6'd75,6'd76,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd62: Enemy_img = 4'd13;
//6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd66,6'd69,6'd70,6'd71,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd62: Enemy_img = 4'd13;
//6'd47,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd69,6'd71,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd61: Enemy_img = 4'd13;
//6'd46,6'd47,6'd49,6'd50,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd64,6'd66,6'd67,6'd68,6'd69,6'd75,6'd76,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd59: Enemy_img = 4'd13;
//6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd73,6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd71,6'd72,6'd76,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd61: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd69,6'd70,6'd76,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd73,6'd74,6'd75,6'd77,6'd78,6'd81: Enemy_img = 4'd14;
//6'd71,6'd72,6'd76,6'd80,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd57,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd55,6'd56,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd75,6'd77,6'd78,6'd79,6'd82: Enemy_img = 4'd14;
//6'd73,6'd74,6'd76,6'd81,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd77,6'd78,6'd79,6'd82,6'd83: Enemy_img = 4'd14;
//6'd75,6'd76,6'd81,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd66,6'd67: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd51,6'd52,6'd56,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd79,6'd80,6'd83,6'd84: Enemy_img = 4'd14;
//6'd76,6'd77,6'd78,6'd82,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd53,6'd54,6'd55,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd56,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd79,6'd80,6'd83,6'd84,6'd86: Enemy_img = 4'd14;
//6'd75,6'd78,6'd82,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd9;
//6'd51,6'd54,6'd55,6'd57: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd56,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd66,6'd74,6'd78,6'd83,6'd84,6'd85,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd9;
//6'd62: Enemy_img = 4'd10;
//6'd52,6'd55: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd56,6'd57,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd65,6'd66,6'd73,6'd78,6'd79,6'd80,6'd81,6'd83,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd64,6'd65: Enemy_img = 4'd9;
//6'd61,6'd62,6'd63: Enemy_img = 4'd10;
//6'd53,6'd57,6'd58: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92: Enemy_img = 4'd14;
//6'd72,6'd82,6'd84,6'd91,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd56,6'd57,6'd58: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd59,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd85,6'd86,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd72,6'd82,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd57,6'd58,6'd60,6'd61,6'd66,6'd67: Enemy_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd59,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd83,6'd86,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd71,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd87,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd88,6'd89,6'd91: Enemy_img = 4'd14;
//6'd71,6'd76,6'd85,6'd86,6'd87,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd9;
//6'd57: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd66,6'd71,6'd76,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd9;
//6'd62: Enemy_img = 4'd10;
//6'd54,6'd57: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd68,6'd69,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd65,6'd66,6'd71,6'd72,6'd73,6'd76,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd64,6'd65: Enemy_img = 4'd9;
//6'd61,6'd62,6'd63: Enemy_img = 4'd10;
//6'd55,6'd58: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85: Enemy_img = 4'd14;
//6'd70,6'd73,6'd76,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd58: Enemy_img = 4'd13;
//6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd59,6'd66,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//6'd70,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd58,6'd60,6'd61,6'd66,6'd67: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd59,6'd62,6'd63,6'd64,6'd65,6'd68,6'd71,6'd72,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd70,6'd73,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd68,6'd71,6'd72,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd70,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd9;
//6'd55: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79: Enemy_img = 4'd14;
//6'd66,6'd70,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd9;
//6'd62: Enemy_img = 4'd10;
//6'd57: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd65,6'd66,6'd71,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd64,6'd65: Enemy_img = 4'd9;
//6'd61,6'd62,6'd63: Enemy_img = 4'd10;
//6'd53,6'd56,6'd57,6'd58: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd72,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd54,6'd59,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd54,6'd55,6'd56,6'd60,6'd61: Enemy_img = 4'd13;
//6'd49,6'd50,6'd53,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76: Enemy_img = 4'd14;
//6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd56,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd50,6'd51,6'd54,6'd55,6'd57,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75: Enemy_img = 4'd14;
//6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd58: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd60,6'd61: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd74: Enemy_img = 4'd14;
//6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd68,6'd69,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd58,6'd59: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd60,6'd62: Enemy_img = 4'd13;
//6'd52,6'd53,6'd57,6'd58,6'd59,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd62: Enemy_img = 4'd13;
//6'd52,6'd58,6'd59,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd56,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd54,6'd55,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd51,6'd52,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73: Enemy_img = 4'd14;
//6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd56,6'd59,6'd60,6'd62: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd55,6'd63,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd62: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd63,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd56,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd53,6'd56,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd59,6'd62: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd73,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd66,6'd67: Enemy_img = 4'd14;
//6'd65,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59: Enemy_img = 4'd14;
//6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd14;
//6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd13;
//6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd13;
//6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd13;
//6'd47: Enemy_img = 4'd14;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd48: Enemy_img = 4'd14;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd46,6'd47,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd47,6'd49,6'd50: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd47,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51: Enemy_img = 4'd14;
//6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51,6'd52: Enemy_img = 4'd14;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51,6'd52: Enemy_img = 4'd14;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51,6'd52,6'd53: Enemy_img = 4'd14;
//6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52,6'd53: Enemy_img = 4'd14;
//6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd13;
//6'd49,6'd50,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53: Enemy_img = 4'd13;
//6'd50,6'd51,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd51,6'd52,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd58,6'd59,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd59,6'd60,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd67: Enemy_img = 4'd13;
//6'd52,6'd53,6'd55,6'd56,6'd57,6'd66,6'd68,6'd69: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd64,6'd65,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd67: Enemy_img = 4'd13;
//6'd50,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd66,6'd68,6'd69: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd64,6'd65,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd68: Enemy_img = 4'd13;
//6'd50,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd61,6'd66,6'd67,6'd69,6'd70: Enemy_img = 4'd14;
//6'd60,6'd62,6'd63,6'd65,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd68: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd58,6'd61,6'd62,6'd69,6'd70: Enemy_img = 4'd14;
//6'd60,6'd63,6'd64,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56: Enemy_img = 4'd13;
//6'd50,6'd51,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd63,6'd70,6'd71: Enemy_img = 4'd14;
//6'd60,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd57,6'd58,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd67,6'd68,6'd69,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd55,6'd57,6'd58,6'd59,6'd62,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd61,6'd63,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd56,6'd58,6'd59,6'd62,6'd64,6'd65,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd48,6'd61,6'd63,6'd66,6'd67,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd13;
//6'd45,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd62,6'd63,6'd66,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd61,6'd64,6'd65,6'd67,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd58: Enemy_img = 4'd13;
//6'd45,6'd46,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd47,6'd48,6'd62,6'd66,6'd67,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd58: Enemy_img = 4'd13;
//6'd43,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd59,6'd60,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd72,6'd73: Enemy_img = 4'd14;
//6'd41,6'd42,6'd47,6'd48,6'd62,6'd66,6'd71,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd58: Enemy_img = 4'd13;
//6'd43,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd59,6'd60,6'd61,6'd63,6'd64,6'd67,6'd68,6'd71,6'd72,6'd73,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd41,6'd42,6'd65,6'd66,6'd70,6'd74,6'd78,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd59: Enemy_img = 4'd13;
//6'd44,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd60,6'd61,6'd63,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd81,6'd82,6'd85,6'd95: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd64,6'd65,6'd69,6'd74,6'd79,6'd80,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd59: Enemy_img = 4'd13;
//6'd44,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd60,6'd61,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd42,6'd43,6'd63,6'd68,6'd74,6'd80,6'd81,6'd84,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd59: Enemy_img = 4'd13;
//6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd65,6'd73,6'd76,6'd77,6'd78,6'd79,6'd85,6'd86,6'd87,6'd88,6'd89,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd42,6'd43,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd82,6'd83,6'd84,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86,6'd87,6'd92: Enemy_img = 4'd14;
//6'd43,6'd44,6'd75,6'd76,6'd77,6'd83,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd79,6'd85,6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd14;
//6'd44,6'd75,6'd78,6'd80,6'd81,6'd84,6'd88,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd52,6'd57,6'd60: Enemy_img = 4'd13;
//6'd47,6'd51,6'd53,6'd54,6'd55,6'd56,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd80,6'd81,6'd87,6'd89,6'd90: Enemy_img = 4'd14;
//6'd45,6'd74,6'd78,6'd79,6'd82,6'd83,6'd85,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd59,6'd60: Enemy_img = 4'd13;
//6'd56,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd74,6'd82,6'd83,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd59,6'd60,6'd61,6'd66,6'd67: Enemy_img = 4'd13;
//6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd83,6'd84,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd80,6'd81,6'd82,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd59,6'd60,6'd61,6'd65: Enemy_img = 4'd13;
//6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd58,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88: Enemy_img = 4'd14;
//6'd73,6'd78,6'd79,6'd80,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd13;
//6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd56,6'd58,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87: Enemy_img = 4'd14;
//6'd67,6'd73,6'd78,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd56,6'd57,6'd60,6'd61,6'd62: Enemy_img = 4'd13;
//6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd55,6'd58,6'd59,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd66,6'd67,6'd73,6'd78,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66: Enemy_img = 4'd9;
//6'd63,6'd64: Enemy_img = 4'd10;
//6'd51,6'd52,6'd55,6'd56: Enemy_img = 4'd13;
//6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd54,6'd57,6'd58,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd73,6'd78,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65: Enemy_img = 4'd10;
//6'd51,6'd54,6'd55,6'd56,6'd58,6'd69: Enemy_img = 4'd13;
//6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd53,6'd57,6'd68,6'd70,6'd71,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd14;
//6'd73,6'd74,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd9;
//6'd63: Enemy_img = 4'd10;
//6'd50,6'd55,6'd56,6'd57,6'd68: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd52,6'd53,6'd54,6'd58,6'd59,6'd66,6'd67,6'd71,6'd72,6'd77,6'd78,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd74,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd57,6'd60,6'd64,6'd66,6'd67: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd55,6'd56,6'd58,6'd59,6'd65,6'd71,6'd72,6'd75,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd69,6'd74,6'd76,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd58,6'd62,6'd71,6'd72,6'd75,6'd76,6'd78,6'd82,6'd83: Enemy_img = 4'd14;
//6'd69,6'd74,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69: Enemy_img = 4'd9;
//6'd55,6'd56,6'd59,6'd60,6'd61: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd71,6'd72,6'd75,6'd76,6'd80,6'd83: Enemy_img = 4'd14;
//6'd74,6'd77,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd67,6'd68: Enemy_img = 4'd9;
//6'd65,6'd66: Enemy_img = 4'd10;
//6'd57,6'd60,6'd61: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd70,6'd71,6'd72,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd74,6'd75,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64: Enemy_img = 4'd9;
//6'd65,6'd66: Enemy_img = 4'd10;
//6'd58,6'd61,6'd71: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd70,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd70: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd67,6'd68,6'd69,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61,6'd62,6'd64,6'd73,6'd74,6'd75,6'd76,6'd81,6'd82: Enemy_img = 4'd14;
//6'd71,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70: Enemy_img = 4'd9;
//6'd60,6'd63,6'd65,6'd66,6'd67: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd64,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82: Enemy_img = 4'd14;
//6'd71,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71: Enemy_img = 4'd9;
//6'd68: Enemy_img = 4'd10;
//6'd60: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67: Enemy_img = 4'd9;
//6'd68,6'd69: Enemy_img = 4'd10;
//6'd61: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd14;
//6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67: Enemy_img = 4'd9;
//6'd61,6'd64: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd68: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd67,6'd68: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd65,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd66,6'd69: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd14;
//6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd13;
//6'd57,6'd58,6'd59,6'd60,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd72: Enemy_img = 4'd13;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd13;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd72,6'd73: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd68,6'd69,6'd70,6'd74,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd70,6'd73: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd68,6'd69,6'd71,6'd74,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd67,6'd68,6'd70,6'd73: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66,6'd69,6'd71,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd70,6'd71,6'd74: Enemy_img = 4'd13;
//6'd69,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd74: Enemy_img = 4'd13;
//6'd63,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd71,6'd75: Enemy_img = 4'd13;
//6'd62,6'd63,6'd67,6'd68,6'd69,6'd70,6'd72,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd72,6'd75: Enemy_img = 4'd13;
//6'd62,6'd63,6'd68,6'd71,6'd73,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd70,6'd72,6'd75: Enemy_img = 4'd13;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd71,6'd73,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd67,6'd70,6'd73,6'd76: Enemy_img = 4'd13;
//6'd61,6'd62,6'd63,6'd66,6'd68,6'd69,6'd71,6'd72,6'd74,6'd77,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd69,6'd70,6'd71,6'd73,6'd76: Enemy_img = 4'd13;
//6'd60,6'd61,6'd62,6'd66,6'd67,6'd68,6'd72,6'd74,6'd77,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd77: Enemy_img = 4'd13;
//6'd59,6'd60,6'd61,6'd66,6'd72,6'd74,6'd75,6'd78: Enemy_img = 4'd14;
//6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd77: Enemy_img = 4'd13;
//6'd58,6'd59,6'd60,6'd66,6'd73,6'd74,6'd75,6'd78: Enemy_img = 4'd14;
//6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63,6'd65: Enemy_img = 4'd13;
//6'd57,6'd58,6'd59,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32: Enemy_img = 4'd13;
//6'd33: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33: Enemy_img = 4'd13;
//6'd34: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36: Enemy_img = 4'd13;
//6'd35,6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37: Enemy_img = 4'd13;
//6'd35,6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd14;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38: Enemy_img = 4'd13;
//6'd36,6'd37,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39: Enemy_img = 4'd13;
//6'd37,6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd43,6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40: Enemy_img = 4'd13;
//6'd38,6'd39,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd44,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd13;
//6'd39,6'd40,6'd42,6'd43,6'd44,6'd60,6'd61: Enemy_img = 4'd14;
//6'd45,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd59: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd60,6'd61: Enemy_img = 4'd14;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd59,6'd60: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd58,6'd61,6'd62,6'd90: Enemy_img = 4'd14;
//6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd60,6'd61: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd59,6'd62,6'd63,6'd89: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd57,6'd58,6'd64,6'd65,6'd66,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd61,6'd62: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd60,6'd63,6'd64,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd65,6'd66,6'd67,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd83,6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd61,6'd62,6'd69,6'd72,6'd73,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88: Enemy_img = 4'd14;
//6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd88: Enemy_img = 4'd14;
//6'd54,6'd62,6'd63,6'd72,6'd73,6'd79,6'd80,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd78,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd62,6'd67,6'd70,6'd75,6'd76,6'd77,6'd79,6'd80,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd44,6'd45,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd57,6'd64,6'd65,6'd68,6'd71,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82,6'd83,6'd86,6'd87: Enemy_img = 4'd14;
//6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd69,6'd70,6'd78,6'd79,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd13;
//6'd45,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd58,6'd61,6'd65,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd83,6'd86,6'd87: Enemy_img = 4'd14;
//6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd67,6'd70,6'd71,6'd81,6'd82,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd45,6'd46,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd73,6'd75,6'd76,6'd77,6'd85,6'd86: Enemy_img = 4'd14;
//6'd57,6'd58,6'd62,6'd66,6'd71,6'd72,6'd74,6'd78,6'd79,6'd80,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd13;
//6'd46,6'd47,6'd51,6'd52,6'd54,6'd55,6'd56,6'd60,6'd61,6'd64,6'd67,6'd68,6'd69,6'd70,6'd71,6'd78,6'd79,6'd82,6'd85,6'd86: Enemy_img = 4'd14;
//6'd58,6'd59,6'd62,6'd63,6'd66,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd55,6'd56,6'd57,6'd60,6'd61,6'd63,6'd64,6'd67,6'd74,6'd75,6'd78,6'd79,6'd82,6'd85,6'd86: Enemy_img = 4'd14;
//6'd59,6'd62,6'd66,6'd68,6'd69,6'd70,6'd73,6'd76,6'd77,6'd80,6'd81,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd58,6'd60,6'd63,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd61,6'd62,6'd65,6'd66,6'd67,6'd73,6'd79,6'd80,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd57,6'd58,6'd59,6'd62,6'd63,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd45,6'd61,6'd65,6'd73,6'd78,6'd79,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd58,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd44,6'd45,6'd59,6'd60,6'd73,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd13;
//6'd43,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd44,6'd45,6'd73,6'd77,6'd78,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd84: Enemy_img = 4'd14;
//6'd45,6'd73,6'd78,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd66: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd83,6'd84: Enemy_img = 4'd14;
//6'd73,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd60,6'd66: Enemy_img = 4'd13;
//6'd41,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd40,6'd74,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd57,6'd60,6'd61,6'd65: Enemy_img = 4'd13;
//6'd42,6'd43,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd78,6'd79,6'd80,6'd84: Enemy_img = 4'd14;
//6'd40,6'd41,6'd67,6'd74,6'd75,6'd76,6'd77,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65: Enemy_img = 4'd13;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd63,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd67,6'd75,6'd76,6'd78,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68: Enemy_img = 4'd9;
//6'd53,6'd54,6'd60,6'd61,6'd62,6'd63,6'd64,6'd70,6'd71: Enemy_img = 4'd13;
//6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd58,6'd59,6'd72,6'd73,6'd74,6'd77,6'd78,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd9;
//6'd65,6'd66: Enemy_img = 4'd10;
//6'd49,6'd50,6'd56,6'd58,6'd61,6'd62,6'd63,6'd70: Enemy_img = 4'd13;
//6'd45,6'd47,6'd48,6'd59,6'd60,6'd69,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd9;
//6'd65,6'd66: Enemy_img = 4'd10;
//6'd55,6'd58,6'd59,6'd70: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd57,6'd60,6'd61,6'd68,6'd69,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd45,6'd71,6'd72,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd9;
//6'd55,6'd58,6'd69: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd59,6'd60,6'd67,6'd68,6'd74,6'd75,6'd80,6'd81,6'd82,6'd83,6'd85: Enemy_img = 4'd14;
//6'd46,6'd71,6'd72,6'd78,6'd79,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72: Enemy_img = 4'd9;
//6'd55,6'd58,6'd61,6'd67,6'd68,6'd75: Enemy_img = 4'd13;
//6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd59,6'd60,6'd74,6'd76,6'd85,6'd86: Enemy_img = 4'd14;
//6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd9;
//6'd57,6'd58,6'd59,6'd63,6'd66,6'd67,6'd74: Enemy_img = 4'd13;
//6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd60,6'd61,6'd62,6'd64,6'd65,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86: Enemy_img = 4'd14;
//6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71: Enemy_img = 4'd10;
//6'd54,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd74: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd56,6'd61,6'd65,6'd73,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd14;
//6'd76,6'd84,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69: Enemy_img = 4'd9;
//6'd70: Enemy_img = 4'd10;
//6'd54,6'd62,6'd63,6'd64,6'd65,6'd73,6'd74: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd72,6'd78,6'd79,6'd80,6'd81,6'd82,6'd87: Enemy_img = 4'd14;
//6'd76,6'd84,6'd85,6'd86,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd75,6'd76: Enemy_img = 4'd9;
//6'd54,6'd59,6'd65,6'd71,6'd72,6'd73: Enemy_img = 4'd13;
//6'd47,6'd48,6'd51,6'd52,6'd53,6'd62,6'd63,6'd64,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87,6'd88,6'd100: Enemy_img = 4'd14;
//6'd84,6'd98,6'd99,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd9;
//6'd60,6'd61,6'd62,6'd66,6'd67,6'd70,6'd71,6'd72: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd64,6'd65,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd83,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74,6'd75: Enemy_img = 4'd10;
//6'd68,6'd71: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd69,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd83,6'd91,6'd92,6'd93,6'd94,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73: Enemy_img = 4'd9;
//6'd74: Enemy_img = 4'd10;
//6'd64,6'd65: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd68,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd83,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd9;
//6'd66,6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd69,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd70,6'd71,6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd76,6'd77,6'd78,6'd79,6'd80,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd82,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd70,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd76,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72,6'd74,6'd77: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd73,6'd75,6'd76,6'd78,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72,6'd74,6'd80: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd73,6'd75,6'd76,6'd77,6'd81,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd70,6'd71,6'd72,6'd81: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd82,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd75,6'd76,6'd77,6'd82: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd78,6'd79,6'd83,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd73,6'd74,6'd83: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd70,6'd76,6'd79,6'd80,6'd84: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd81,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd79,6'd86,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd86: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd69,6'd70,6'd71,6'd72,6'd73,6'd80,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd77,6'd83,6'd87: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd71,6'd72,6'd73,6'd74,6'd76,6'd81,6'd84,6'd88,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd77,6'd83,6'd84,6'd88: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd79,6'd80,6'd81,6'd82,6'd85,6'd89,6'd92,6'd93: Enemy_img = 4'd14;
//6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd82,6'd84,6'd85,6'd89: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd79,6'd80,6'd81,6'd83,6'd86,6'd90: Enemy_img = 4'd14;
//6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd83,6'd85,6'd86,6'd90: Enemy_img = 4'd13;
//6'd44,6'd75,6'd76,6'd81,6'd82,6'd84,6'd87,6'd91: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd13;
//6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd85,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd13;
//6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd13;
//6'd75,6'd76,6'd79,6'd80,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd13;
//6'd74,6'd75,6'd76,6'd80,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd13;
//6'd74,6'd75,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd13;
//6'd74,6'd75,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77: Enemy_img = 4'd13;
//6'd73,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd13;
//6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd14;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81: Enemy_img = 4'd14;
//6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81: Enemy_img = 4'd14;
//6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80: Enemy_img = 4'd14;
//6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd14;
//6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd73,6'd74,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56,6'd72,6'd73,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd69,6'd70,6'd71,6'd72,6'd73,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd80,6'd81: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd13;
//6'd23,6'd24,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd80,6'd81: Enemy_img = 4'd14;
//6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd23,6'd24,6'd53,6'd54,6'd55: Enemy_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd51,6'd52,6'd56,6'd57,6'd77,6'd81: Enemy_img = 4'd14;
//6'd60,6'd75,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd53,6'd54,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd51,6'd52,6'd58,6'd59,6'd60,6'd65,6'd73,6'd74,6'd76,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29: Enemy_img = 4'd13;
//6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd59,6'd60,6'd61,6'd63,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd55,6'd56,6'd57,6'd58,6'd62,6'd64,6'd65,6'd70,6'd73,6'd76,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd27,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd56,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd38,6'd39,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd62,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd13;
//6'd30,6'd31,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd62,6'd68,6'd69,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd63,6'd64,6'd65,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd57,6'd58,6'd59,6'd62,6'd66,6'd67,6'd75,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd51,6'd55,6'd57,6'd60,6'd61,6'd64,6'd68,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd14;
//6'd50,6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd63,6'd65,6'd66,6'd70,6'd75,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41: Enemy_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd53,6'd54,6'd57,6'd60,6'd61,6'd63,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd78,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd51,6'd52,6'd55,6'd56,6'd58,6'd59,6'd64,6'd65,6'd70,6'd75,6'd76,6'd77,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43: Enemy_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd55,6'd56,6'd57,6'd58,6'd61,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd83: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd59,6'd60,6'd63,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd51,6'd57,6'd58,6'd60,6'd61,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd59,6'd63,6'd71,6'd80,6'd81,6'd82,6'd83,6'd84,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd57,6'd59,6'd72,6'd76,6'd80,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55,6'd56,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd81,6'd82,6'd83,6'd84,6'd85,6'd101: Enemy_img = 4'd14;
//6'd59,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd100,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd66: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd57,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd100,6'd101: Enemy_img = 4'd14;
//6'd58,6'd75,6'd99,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd65: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd86,6'd87,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd76,6'd83,6'd84,6'd85,6'd98,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd65: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd79,6'd80,6'd86,6'd87,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd67,6'd77,6'd78,6'd81,6'd85,6'd88,6'd97,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd9;
//6'd57,6'd65,6'd71: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd70,6'd74,6'd75,6'd76,6'd82,6'd83,6'd84,6'd89,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd67,6'd79,6'd86,6'd87,6'd88,6'd95,6'd96,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd9;
//6'd60,6'd65,6'd71: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd61,6'd62,6'd63,6'd64,6'd70,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd88,6'd89,6'd90,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd73,6'd86,6'd87,6'd93,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd9;
//6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd71,6'd76: Enemy_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd70,6'd75,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd44,6'd73,6'd86,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd9;
//6'd66,6'd67: Enemy_img = 4'd10;
//6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd71,6'd76: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd69,6'd70,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd44,6'd45,6'd78,6'd86,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd72,6'd73: Enemy_img = 4'd9;
//6'd67: Enemy_img = 4'd10;
//6'd61,6'd62,6'd63,6'd70: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd69,6'd76,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd78,6'd79,6'd86,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd78,6'd79: Enemy_img = 4'd9;
//6'd72,6'd73: Enemy_img = 4'd10;
//6'd56,6'd69,6'd70,6'd76: Enemy_img = 4'd13;
//6'd43,6'd44,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd75,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd45,6'd46,6'd86,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd78,6'd79: Enemy_img = 4'd9;
//6'd72,6'd73: Enemy_img = 4'd10;
//6'd54,6'd55,6'd58,6'd60,6'd61,6'd68,6'd69,6'd76: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd59,6'd62,6'd75,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd86,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd9;
//6'd78,6'd79: Enemy_img = 4'd10;
//6'd42,6'd43,6'd44,6'd57,6'd58,6'd60,6'd61,6'd63,6'd66,6'd67,6'd74,6'd75: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd59,6'd62,6'd64,6'd68,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd77: Enemy_img = 4'd9;
//6'd78: Enemy_img = 4'd10;
//6'd45,6'd46,6'd52,6'd53,6'd58,6'd60,6'd61,6'd62,6'd66,6'd67,6'd68,6'd74,6'd75: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd47,6'd49,6'd50,6'd51,6'd54,6'd56,6'd57,6'd63,6'd64,6'd65,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77: Enemy_img = 4'd9;
//6'd78: Enemy_img = 4'd10;
//6'd47,6'd48,6'd51,6'd52,6'd58,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72: Enemy_img = 4'd13;
//6'd45,6'd46,6'd50,6'd54,6'd55,6'd56,6'd57,6'd60,6'd65,6'd73,6'd74,6'd80,6'd81,6'd82,6'd83,6'd84,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77: Enemy_img = 4'd9;
//6'd58,6'd61,6'd62,6'd73,6'd79,6'd80: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd79,6'd80,6'd82,6'd86,6'd87: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd72,6'd73,6'd74,6'd78,6'd81,6'd83,6'd88,6'd89,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd62,6'd63,6'd64,6'd65,6'd69,6'd70,6'd71,6'd76,6'd77,6'd80,6'd82,6'd88,6'd89: Enemy_img = 4'd13;
//6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd66,6'd67,6'd68,6'd75,6'd78,6'd79,6'd81,6'd83,6'd90,6'd91,6'd92,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd49,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd72,6'd73,6'd76,6'd77,6'd80,6'd84,6'd90,6'd91,6'd92: Enemy_img = 4'd13;
//6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd78,6'd79,6'd81,6'd85,6'd86,6'd93,6'd94,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd74,6'd76,6'd77,6'd78,6'd79,6'd83,6'd89,6'd92,6'd93,6'd94: Enemy_img = 4'd13;
//6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd80,6'd84,6'd85,6'd86,6'd87,6'd88,6'd95,6'd96: Enemy_img = 4'd14;
//6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd81,6'd82,6'd87,6'd88,6'd89,6'd95,6'd96,6'd97: Enemy_img = 4'd13;
//6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd79,6'd83,6'd84,6'd85,6'd86,6'd92,6'd98,6'd99: Enemy_img = 4'd14;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd77,6'd80,6'd81,6'd84,6'd85,6'd86,6'd91,6'd97,6'd98,6'd99: Enemy_img = 4'd13;
//6'd53,6'd54,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd78,6'd82,6'd83,6'd87,6'd88,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd92,6'd93,6'd94: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd80,6'd81,6'd89,6'd90,6'd91,6'd95,6'd96: Enemy_img = 4'd14;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd86,6'd90,6'd91,6'd95,6'd96: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd79,6'd80,6'd81,6'd85,6'd89,6'd92,6'd93,6'd94,6'd97,6'd98: Enemy_img = 4'd14;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84,6'd86,6'd92,6'd93: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd88,6'd89,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd91,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd89,6'd90,6'd92,6'd93,6'd94: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd85,6'd88,6'd91,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd92,6'd93,6'd94: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd89,6'd92,6'd93: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd85,6'd86,6'd87,6'd90,6'd91,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd89,6'd90: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd85,6'd86,6'd87,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd86,6'd87,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd89,6'd90: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd86,6'd87,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd89,6'd90: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd86,6'd87,6'd91,6'd92: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88,6'd89: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd86,6'd87,6'd90,6'd91: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd88: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd86,6'd87,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd86,6'd87: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd86: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72: Enemy_img = 4'd14;
//6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72: Enemy_img = 4'd14;
//6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd14;
//6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70: Enemy_img = 4'd14;
//6'd68,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd67,6'd68,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd67,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd70,6'd74,6'd75: Enemy_img = 4'd14;
//6'd66,6'd67,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd14;
//6'd66,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd65,6'd66,6'd67,6'd68,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd69,6'd76: Enemy_img = 4'd14;
//6'd64,6'd65,6'd68,6'd70,6'd71,6'd74,6'd75,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd72,6'd73: Enemy_img = 4'd14;
//6'd63,6'd64,6'd68,6'd69,6'd76,6'd77,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd73,6'd74,6'd75,6'd99: Enemy_img = 4'd14;
//6'd62,6'd63,6'd66,6'd67,6'd70,6'd71,6'd72,6'd98,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd99: Enemy_img = 4'd14;
//6'd61,6'd62,6'd64,6'd65,6'd69,6'd72,6'd77,6'd98,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd63,6'd69,6'd72,6'd77,6'd97,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd59,6'd60,6'd61,6'd69,6'd72,6'd77,6'd97,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd66,6'd67,6'd68,6'd69,6'd72,6'd77,6'd96,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd78,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd61,6'd66,6'd72,6'd77,6'd79,6'd80,6'd81,6'd82,6'd96,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd60,6'd67,6'd68,6'd69,6'd70,6'd71,6'd80,6'd81,6'd82,6'd83,6'd84,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd56,6'd57,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd95,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd55,6'd56,6'd59,6'd65,6'd67,6'd79,6'd94,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd89,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd54,6'd55,6'd60,6'd64,6'd68,6'd79,6'd84,6'd88,6'd93,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82,6'd86,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd60,6'd64,6'd69,6'd75,6'd76,6'd77,6'd78,6'd79,6'd83,6'd85,6'd87,6'd88,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd56,6'd57,6'd58,6'd59,6'd62,6'd65,6'd66,6'd67,6'd68,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd88,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd52,6'd53,6'd55,6'd61,6'd63,6'd70,6'd71,6'd75,6'd82,6'd86,6'd87,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd59,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd76,6'd77,6'd78,6'd79,6'd80,6'd83,6'd84,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd48,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd61,6'd63,6'd72,6'd73,6'd74,6'd75,6'd81,6'd87,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd60,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd82,6'd83,6'd84,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd55,6'd57,6'd62,6'd76,6'd77,6'd78,6'd79,6'd80,6'd87,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd60,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd55,6'd57,6'd58,6'd59,6'd62,6'd88,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd88,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd72,6'd78: Enemy_img = 4'd13;
//6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd70,6'd71,6'd76,6'd77,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd59,6'd89,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd72,6'd78: Enemy_img = 4'd13;
//6'd58,6'd60,6'd62,6'd63,6'd64,6'd65,6'd71,6'd77,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd68,6'd69,6'd74,6'd75,6'd80,6'd81,6'd89,6'd106,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd76,6'd82: Enemy_img = 4'd9;
//6'd67,6'd73,6'd79: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd62,6'd63,6'd64,6'd65,6'd66,6'd72,6'd78,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd69,6'd75,6'd81,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd75,6'd76,6'd81,6'd82: Enemy_img = 4'd9;
//6'd67,6'd73,6'd79: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd72,6'd78,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd59,6'd68,6'd71,6'd74,6'd77,6'd80,6'd83,6'd89,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd69,6'd75,6'd81: Enemy_img = 4'd9;
//6'd70,6'd76,6'd82: Enemy_img = 4'd10;
//6'd67,6'd73,6'd79: Enemy_img = 4'd13;
//default: Enemy_img = 4'd14;
//endcase
//end
//6'd64: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd59,6'd68,6'd71,6'd74,6'd77,6'd80,6'd83,6'd89,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd69,6'd70,6'd75,6'd76,6'd81,6'd82: Enemy_img = 4'd10;
//default: Enemy_img = 4'd13;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd72,6'd78,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd75,6'd81: Enemy_img = 4'd9;
//6'd70,6'd76,6'd82: Enemy_img = 4'd10;
//6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd78,6'd79,6'd84,6'd85,6'd87: Enemy_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd86,6'd88: Enemy_img = 4'd14;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd75,6'd76,6'd81,6'd82: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd78,6'd79,6'd84,6'd85,6'd87,6'd90,6'd95: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd62,6'd86,6'd88,6'd91,6'd92,6'd93,6'd94,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd74,6'd75,6'd80,6'd81: Enemy_img = 4'd9;
//6'd60,6'd63,6'd64,6'd65,6'd66,6'd85,6'd89,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd71,6'd72,6'd77,6'd78,6'd83,6'd84,6'd86,6'd87,6'd90,6'd91,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd70,6'd71,6'd72,6'd76,6'd77,6'd78,6'd82,6'd83,6'd85,6'd86,6'd89: Enemy_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd84,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd81,6'd82,6'd83,6'd88,6'd91,6'd92,6'd93,6'd94,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd66,6'd69,6'd76,6'd77,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86,6'd89,6'd90,6'd96,6'd104,6'd105: Enemy_img = 4'd14;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd62,6'd65,6'd71,6'd82,6'd83,6'd84,6'd85,6'd88,6'd90,6'd91,6'd92,6'd93,6'd95,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd81,6'd86,6'd89,6'd96,6'd97,6'd98,6'd99,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd76,6'd77,6'd78,6'd79,6'd80,6'd83,6'd84,6'd87,6'd90,6'd91,6'd93,6'd97,6'd98,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd64,6'd70,6'd71,6'd82,6'd85,6'd88,6'd89,6'd92,6'd95,6'd96,6'd99,6'd103,6'd104: Enemy_img = 4'd14;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd63,6'd66,6'd67,6'd68,6'd72,6'd73,6'd75,6'd84,6'd89,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd65,6'd69,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd85,6'd87,6'd88,6'd92,6'd99,6'd103,6'd104: Enemy_img = 4'd14;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd66,6'd67,6'd70,6'd71,6'd82,6'd86,6'd91,6'd92,6'd94,6'd95,6'd100,6'd101: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd65,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd87,6'd88,6'd89,6'd90,6'd96,6'd97,6'd98,6'd99,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd64,6'd69,6'd83,6'd85,6'd95,6'd97,6'd98: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd96,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd64,6'd68,6'd84,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd93,6'd94,6'd95,6'd96,6'd102,6'd103: Enemy_img = 4'd14;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd65,6'd67,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd94,6'd95,6'd96,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd66,6'd98,6'd99,6'd100: Enemy_img = 4'd13;
//6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd95,6'd96,6'd97,6'd101,6'd102: Enemy_img = 4'd14;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd98,6'd99,6'd100: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd96,6'd97,6'd101,6'd102: Enemy_img = 4'd14;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd99: Enemy_img = 4'd13;
//6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd99: Enemy_img = 4'd13;
//6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd97,6'd98,6'd100,6'd101: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd76,6'd77,6'd99: Enemy_img = 4'd14;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd99: Enemy_img = 4'd14;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_3 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd14;
//6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd88: Enemy_img = 4'd14;
//6'd57,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd88,6'd89: Enemy_img = 4'd14;
//6'd57,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd57,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd87,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd61,6'd62,6'd63,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd57,6'd60,6'd87,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd57,6'd60,6'd61,6'd87,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd64,6'd65,6'd66,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd57,6'd61,6'd62,6'd63,6'd87,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd56,6'd57,6'd63,6'd64,6'd87,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd56,6'd62,6'd67,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd64,6'd65,6'd66,6'd67,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59,6'd61,6'd68,6'd86,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd69,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd56,6'd59,6'd60,6'd62,6'd63,6'd64,6'd69,6'd74,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd55,6'd56,6'd59,6'd61,6'd64,6'd69,6'd70,6'd72,6'd73,6'd81,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd60,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd55,6'd58,6'd61,6'd65,6'd70,6'd71,6'd72,6'd77,6'd78,6'd81,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd59,6'd60,6'd61,6'd63,6'd64,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd55,6'd57,6'd62,6'd65,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd78,6'd79,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd100,6'd101: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd73,6'd77,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd101: Enemy_img = 4'd13;
//6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd93,6'd94,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd54,6'd55,6'd60,6'd61,6'd66,6'd72,6'd73,6'd76,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd98,6'd99,6'd100: Enemy_img = 4'd13;
//6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd96,6'd97: Enemy_img = 4'd14;
//6'd53,6'd54,6'd60,6'd70,6'd71,6'd76,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd96,6'd97: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd86,6'd87,6'd88,6'd89,6'd90,6'd93,6'd94,6'd95,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd53,6'd54,6'd59,6'd60,6'd61,6'd70,6'd75,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93,6'd94,6'd95: Enemy_img = 4'd13;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd91,6'd92,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92,6'd93,6'd99,6'd100: Enemy_img = 4'd13;
//6'd55,6'd57,6'd58,6'd59,6'd61,6'd62,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88,6'd89,6'd90,6'd96,6'd97,6'd98,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd50,6'd56,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89,6'd90,6'd96,6'd97,6'd98: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88,6'd95,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd9;
//6'd75,6'd93,6'd95,6'd96,6'd99,6'd100,6'd101: Enemy_img = 4'd13;
//6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd91,6'd92,6'd97,6'd98,6'd102,6'd103: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd55,6'd59,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd9;
//6'd76,6'd92,6'd93,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd13;
//6'd48,6'd49,6'd52,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd75,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90,6'd91,6'd95,6'd96,6'd102,6'd103: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd56,6'd59,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd9;
//6'd80: Enemy_img = 4'd10;
//6'd69,6'd77,6'd85,6'd88,6'd91,6'd96,6'd99,6'd100,6'd101: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd75,6'd76,6'd82,6'd83,6'd84,6'd86,6'd89,6'd90,6'd92,6'd93,6'd95,6'd97,6'd98,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd43,6'd44,6'd50,6'd51,6'd57,6'd59,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd9;
//6'd79,6'd80: Enemy_img = 4'd10;
//6'd48,6'd70,6'd77,6'd82,6'd83,6'd84,6'd86,6'd88,6'd92,6'd93,6'd94,6'd97,6'd100,6'd101: Enemy_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd76,6'd85,6'd89,6'd90,6'd91,6'd95,6'd96,6'd98,6'd99,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd50,6'd51,6'd58,6'd59,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74,6'd80: Enemy_img = 4'd9;
//6'd81: Enemy_img = 4'd10;
//6'd46,6'd47,6'd71,6'd77,6'd78,6'd83,6'd84,6'd88,6'd90,6'd91,6'd92,6'd93,6'd96,6'd97,6'd98,6'd100,6'd101: Enemy_img = 4'd13;
//6'd44,6'd45,6'd51,6'd56,6'd57,6'd61,6'd62,6'd63,6'd69,6'd70,6'd76,6'd85,6'd86,6'd89,6'd95,6'd99,6'd102,6'd103: Enemy_img = 4'd14;
//6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd59,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd80,6'd81: Enemy_img = 4'd9;
//6'd74,6'd75: Enemy_img = 4'd10;
//6'd45,6'd64,6'd71,6'd77,6'd78,6'd84,6'd85,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd13;
//6'd46,6'd47,6'd51,6'd55,6'd57,6'd58,6'd61,6'd62,6'd63,6'd70,6'd83,6'd86,6'd89,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd49,6'd50,6'd52,6'd53,6'd54,6'd56,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69,6'd80: Enemy_img = 4'd9;
//6'd74,6'd75: Enemy_img = 4'd10;
//6'd65,6'd72,6'd77,6'd78,6'd82,6'd88,6'd90,6'd91,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd45,6'd50,6'd51,6'd54,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd71,6'd83,6'd84,6'd85,6'd86,6'd89,6'd92,6'd97,6'd103,6'd104: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd52,6'd53,6'd55,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd74,6'd75: Enemy_img = 4'd9;
//6'd69: Enemy_img = 4'd10;
//6'd66,6'd72,6'd82,6'd83,6'd84,6'd85,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd71,6'd77,6'd78,6'd86,6'd88,6'd89,6'd97,6'd103,6'd104: Enemy_img = 4'd14;
//6'd45,6'd46,6'd48,6'd49,6'd53,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd9;
//6'd68,6'd69: Enemy_img = 4'd10;
//6'd66,6'd72,6'd77,6'd78,6'd82,6'd83,6'd84,6'd85,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd61,6'd62,6'd63,6'd64,6'd65,6'd80,6'd81,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98,6'd103,6'd104: Enemy_img = 4'd14;
//6'd47,6'd48,6'd52,6'd53,6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70: Enemy_img = 4'd9;
//6'd66,6'd67,6'd76,6'd84,6'd85,6'd100,6'd101,6'd102: Enemy_img = 4'd13;
//6'd48,6'd49,6'd51,6'd52,6'd53,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd72,6'd77,6'd78,6'd79,6'd83,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd95,6'd96,6'd97,6'd98,6'd99,6'd103,6'd104: Enemy_img = 4'd14;
//6'd46,6'd47,6'd50,6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70: Enemy_img = 4'd9;
//6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd75,6'd76,6'd80,6'd81,6'd87,6'd101,6'd102: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd51,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd71,6'd77,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91,6'd98,6'd99,6'd100,6'd103,6'd104: Enemy_img = 4'd14;
//6'd45,6'd46,6'd50,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd71,6'd72,6'd73,6'd74,6'd78,6'd79,6'd84,6'd87,6'd102: Enemy_img = 4'd13;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83,6'd88,6'd89,6'd90,6'd99,6'd100,6'd101,6'd103,6'd104: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd63,6'd64,6'd65,6'd66,6'd71,6'd72,6'd73,6'd77,6'd86: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd62,6'd67,6'd70,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd68,6'd69,6'd75,6'd77: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd59,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd62,6'd66,6'd70,6'd71,6'd74: Enemy_img = 4'd13;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57,6'd60,6'd61,6'd64,6'd65,6'd67,6'd68,6'd69,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd103,6'd104: Enemy_img = 4'd14;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd64,6'd68,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd66,6'd67,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd104: Enemy_img = 4'd14;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd63,6'd65,6'd69,6'd72: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd68,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd37,6'd38: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd66,6'd72: Enemy_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd62,6'd67,6'd71: Enemy_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd34: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd68,6'd69,6'd71: Enemy_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd62,6'd70: Enemy_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd62: Enemy_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd36,6'd37,6'd38,6'd39,6'd40,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd62: Enemy_img = 4'd13;
//6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30: Enemy_img = 4'd13;
//6'd26,6'd27,6'd31,6'd32,6'd33,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd28: Enemy_img = 4'd13;
//6'd24,6'd25,6'd29,6'd30,6'd55,6'd56,6'd57,6'd58,6'd77,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd57,6'd58,6'd59: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd13;
//6'd54,6'd58,6'd59,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd13;
//6'd55,6'd56,6'd57,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd58,6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83: Enemy_img = 4'd14;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//2'd4: begin
//case(angle)
//// Enemy_type_4 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd86: Enemy_img = 4'd14;
//6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd6;
//6'd52,6'd53,6'd86: Enemy_img = 4'd14;
//6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd57: Enemy_img = 4'd6;
//6'd54,6'd85,6'd86: Enemy_img = 4'd14;
//6'd52,6'd53,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd57,6'd58,6'd59,6'd83: Enemy_img = 4'd6;
//6'd51,6'd52,6'd54,6'd86: Enemy_img = 4'd14;
//6'd53,6'd55,6'd85,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd58,6'd59,6'd60,6'd61,6'd81,6'd82: Enemy_img = 4'd6;
//6'd51,6'd52,6'd54,6'd55,6'd84: Enemy_img = 4'd14;
//6'd53,6'd56,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd59,6'd60,6'd61,6'd62,6'd63,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd55,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd59,6'd60,6'd81: Enemy_img = 4'd7;
//6'd50,6'd52,6'd53,6'd55,6'd56,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd51,6'd54,6'd57,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd60,6'd61,6'd80,6'd81: Enemy_img = 4'd7;
//6'd49,6'd50,6'd52,6'd53,6'd55,6'd56,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd51,6'd54,6'd57,6'd58,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd47,6'd60,6'd61,6'd62,6'd63,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd49,6'd50,6'd52,6'd53,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd25,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd46,6'd61,6'd62,6'd63,6'd64,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd25,6'd51,6'd52,6'd58,6'd59,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd45,6'd46,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd25,6'd48,6'd55,6'd56,6'd57,6'd58,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd24,6'd26,6'd49,6'd50,6'd53,6'd54,6'd59,6'd60,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd6;
//6'd44,6'd45,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd25,6'd51,6'd52,6'd57,6'd58,6'd59,6'd80,6'd82,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd24,6'd26,6'd47,6'd48,6'd55,6'd56,6'd60,6'd61,6'd81,6'd83,6'd84,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd6;
//6'd29,6'd43,6'd44,6'd45,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd24,6'd25,6'd26,6'd49,6'd51,6'd52,6'd53,6'd59,6'd60,6'd79,6'd80,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd23,6'd27,6'd50,6'd54,6'd57,6'd58,6'd61,6'd62,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd41,6'd42,6'd43,6'd44,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd24,6'd25,6'd26,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd55,6'd56,6'd61,6'd78,6'd79,6'd80,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd23,6'd27,6'd50,6'd54,6'd59,6'd60,6'd62,6'd63,6'd81,6'd82,6'd85,6'd86,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd83,6'd84: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33,6'd39,6'd40,6'd41,6'd42,6'd43,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd45,6'd46,6'd47,6'd48,6'd49,6'd55,6'd56,6'd57,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd22,6'd28,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd61,6'd62,6'd63,6'd64,6'd77,6'd78,6'd79,6'd80,6'd81,6'd86,6'd87,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd67,6'd68,6'd69,6'd70,6'd71,6'd82,6'd83: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd75,6'd76,6'd77,6'd78,6'd89,6'd90: Enemy_img = 4'd14;
//6'd22,6'd28,6'd50,6'd58,6'd63,6'd64,6'd65,6'd79,6'd80,6'd87,6'd88,6'd91,6'd92,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85,6'd86: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd68,6'd69,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54,6'd55,6'd61,6'd62,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd22,6'd29,6'd42,6'd46,6'd47,6'd48,6'd49,6'd50,6'd56,6'd57,6'd58,6'd59,6'd60,6'd65,6'd66,6'd78,6'd79,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd82,6'd83: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd40,6'd41,6'd42,6'd44,6'd45,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd61,6'd62,6'd64,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd89,6'd91,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd21,6'd30,6'd43,6'd46,6'd50,6'd56,6'd60,6'd63,6'd70,6'd79,6'd80,6'd87,6'd88,6'd90,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd47,6'd48,6'd49,6'd57,6'd58,6'd59,6'd64,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd88,6'd89,6'd91,6'd92: Enemy_img = 4'd14;
//6'd21,6'd31,6'd43,6'd46,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd65,6'd67,6'd68,6'd70,6'd80,6'd81,6'd86,6'd87,6'd90,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83: Enemy_img = 4'd6;
//6'd84,6'd85: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd38,6'd39,6'd40,6'd41,6'd42,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd63,6'd64,6'd67,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd89,6'd93,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd21,6'd35,6'd36,6'd37,6'd43,6'd44,6'd45,6'd46,6'd50,6'd62,6'd65,6'd68,6'd69,6'd71,6'd79,6'd80,6'd87,6'd88,6'd90,6'd91,6'd92,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82: Enemy_img = 4'd6;
//6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd60,6'd61,6'd66,6'd67,6'd68,6'd73,6'd74,6'd75,6'd76,6'd77,6'd90,6'd91,6'd93,6'd94,6'd98,6'd99: Enemy_img = 4'd14;
//6'd20,6'd37,6'd38,6'd46,6'd50,6'd62,6'd63,6'd64,6'd69,6'd70,6'd72,6'd78,6'd79,6'd88,6'd89,6'd92,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81: Enemy_img = 4'd6;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd74,6'd91,6'd93: Enemy_img = 4'd14;
//6'd20,6'd38,6'd46,6'd50,6'd64,6'd70,6'd71,6'd73,6'd75,6'd76,6'd77,6'd78,6'd89,6'd90,6'd92,6'd94,6'd95,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82: Enemy_img = 4'd6;
//6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd41,6'd43,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd65,6'd69,6'd70,6'd76,6'd77,6'd90,6'd91: Enemy_img = 4'd14;
//6'd20,6'd38,6'd44,6'd45,6'd46,6'd50,6'd63,6'd66,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75,6'd78,6'd79,6'd88,6'd89,6'd92,6'd93,6'd96,6'd97,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83: Enemy_img = 4'd6;
//6'd84,6'd85: Enemy_img = 4'd7;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd78,6'd89,6'd90,6'd91,6'd94,6'd95,6'd97: Enemy_img = 4'd14;
//6'd19,6'd63,6'd68,6'd72,6'd73,6'd76,6'd77,6'd79,6'd80,6'd87,6'd88,6'd92,6'd96,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd64,6'd65,6'd66,6'd67,6'd72,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd19,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd6;
//6'd83: Enemy_img = 4'd7;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd74,6'd88,6'd89,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd18,6'd71,6'd73,6'd75,6'd76,6'd77,6'd80,6'd81,6'd86,6'd87,6'd90,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd28,6'd38,6'd62,6'd80,6'd81,6'd82,6'd85,6'd90,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//default: Enemy_img = 4'd14;
//6'd17,6'd18,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd77,6'd78,6'd79,6'd86,6'd87,6'd89,6'd100,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd28,6'd37,6'd46,6'd47,6'd48,6'd62,6'd82,6'd85,6'd89,6'd95,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd83: Enemy_img = 4'd6;
//6'd84: Enemy_img = 4'd7;
//default: Enemy_img = 4'd14;
//6'd16,6'd17,6'd67,6'd70,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd82,6'd85,6'd95: Enemy_img = 4'd7;
//6'd46,6'd47: Enemy_img = 4'd9;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd89,6'd90,6'd91,6'd92,6'd93,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd87,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd58: Enemy_img = 4'd2;
//6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd75,6'd76,6'd77,6'd84,6'd85,6'd96: Enemy_img = 4'd6;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd86,6'd94,6'd95: Enemy_img = 4'd7;
//6'd45,6'd46: Enemy_img = 4'd9;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd60,6'd61,6'd62,6'd89,6'd90,6'd91,6'd92,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd88,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd57: Enemy_img = 4'd2;
//6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76,6'd85,6'd86,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd20,6'd25,6'd26,6'd31,6'd32,6'd65,6'd66,6'd71,6'd72,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd93,6'd94: Enemy_img = 4'd7;
//6'd46: Enemy_img = 4'd9;
//6'd45: Enemy_img = 4'd10;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd56: Enemy_img = 4'd2;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd35,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd87,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd66,6'd67,6'd68,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd92,6'd96: Enemy_img = 4'd7;
//6'd45,6'd46: Enemy_img = 4'd10;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd98,6'd99,6'd100,6'd101,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd102,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd56: Enemy_img = 4'd2;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd35,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd87,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd66,6'd67,6'd68,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd90,6'd96: Enemy_img = 4'd7;
//6'd46: Enemy_img = 4'd9;
//6'd45: Enemy_img = 4'd10;
//6'd48: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd57: Enemy_img = 4'd2;
//6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd76,6'd85,6'd86,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd20,6'd25,6'd26,6'd31,6'd32,6'd65,6'd66,6'd71,6'd72,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd93,6'd94: Enemy_img = 4'd7;
//6'd45,6'd46: Enemy_img = 4'd9;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd48,6'd49,6'd50,6'd55,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd37,6'd43,6'd54,6'd63,6'd99,6'd100,6'd101,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd58: Enemy_img = 4'd2;
//6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd75,6'd76,6'd77,6'd84,6'd85,6'd96: Enemy_img = 4'd6;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd86,6'd94,6'd95: Enemy_img = 4'd7;
//6'd45: Enemy_img = 4'd9;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd55,6'd56: Enemy_img = 4'd14;
//6'd37,6'd46,6'd51,6'd60,6'd61,6'd62,6'd89,6'd90,6'd91,6'd101,6'd103,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd82,6'd85,6'd95: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd49,6'd50,6'd52,6'd55,6'd56,6'd57,6'd60,6'd61: Enemy_img = 4'd14;
//6'd35,6'd38,6'd39,6'd40,6'd41,6'd46,6'd47,6'd51,6'd62,6'd64,6'd66,6'd89,6'd93,6'd97,6'd98,6'd99,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83: Enemy_img = 4'd6;
//6'd84: Enemy_img = 4'd7;
//6'd39,6'd40,6'd49,6'd50,6'd57,6'd59,6'd60: Enemy_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd61,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd91,6'd92,6'd93,6'd94,6'd97,6'd98,6'd99,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd40,6'd42,6'd43,6'd44,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd57,6'd59,6'd60: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd41,6'd45,6'd46,6'd47,6'd48,6'd51,6'd56,6'd58,6'd61,6'd63,6'd64,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76,6'd88,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd6;
//6'd83: Enemy_img = 4'd7;
//6'd40,6'd42,6'd43,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd18,6'd19,6'd20,6'd39,6'd41,6'd44,6'd49,6'd50,6'd51,6'd52,6'd56,6'd57,6'd58,6'd59,6'd60,6'd64,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd88,6'd89,6'd92,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd42,6'd55,6'd56,6'd58,6'd59: Enemy_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd43,6'd53,6'd54,6'd57,6'd60,6'd64,6'd65,6'd66,6'd68,6'd70,6'd71,6'd72,6'd88,6'd89,6'd90,6'd94,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83: Enemy_img = 4'd6;
//6'd84,6'd85: Enemy_img = 4'd7;
//6'd41,6'd56,6'd58: Enemy_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd42,6'd45,6'd46,6'd47,6'd48,6'd55,6'd57,6'd59,6'd62,6'd70,6'd71,6'd78,6'd89,6'd90,6'd91,6'd94,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82: Enemy_img = 4'd6;
//6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd58: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd56,6'd57,6'd59,6'd62,6'd65,6'd66,6'd67,6'd68,6'd70,6'd76,6'd77,6'd90,6'd91,6'd96,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81: Enemy_img = 4'd6;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd98,6'd99: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd38,6'd39,6'd43,6'd44,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76,6'd91,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82: Enemy_img = 4'd6;
//6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd98,6'd99: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd34,6'd35,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd73,6'd74,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83: Enemy_img = 4'd6;
//6'd84,6'd85: Enemy_img = 4'd7;
//6'd97,6'd98,6'd99: Enemy_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd30,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd53,6'd54,6'd55,6'd56,6'd57,6'd64,6'd71,6'd72,6'd73,6'd74,6'd79,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd82,6'd83: Enemy_img = 4'd7;
//6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd64,6'd71,6'd72,6'd76,6'd77,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85,6'd86: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd68,6'd69,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd72,6'd74,6'd75,6'd76,6'd77,6'd90,6'd91,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd67,6'd68,6'd69,6'd70,6'd71,6'd82,6'd83: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd75,6'd76,6'd77,6'd78,6'd89,6'd90,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd83,6'd84: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33,6'd39,6'd40,6'd41,6'd42,6'd43,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd58,6'd77,6'd78,6'd79,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd41,6'd42,6'd43,6'd44,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd61,6'd78,6'd79,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd6;
//6'd29,6'd43,6'd44,6'd45,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd49,6'd50,6'd51,6'd59,6'd60,6'd79,6'd81,6'd86,6'd87,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd6;
//6'd44,6'd45,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd24,6'd25,6'd51,6'd52,6'd57,6'd58,6'd59,6'd81,6'd82,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd45,6'd46,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd24,6'd25,6'd48,6'd55,6'd57,6'd58,6'd81,6'd82,6'd83,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd46,6'd61,6'd62,6'd63,6'd64,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd82,6'd83,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd47,6'd60,6'd61,6'd62,6'd63,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd60,6'd61,6'd80,6'd81: Enemy_img = 4'd7;
//6'd49,6'd50,6'd54,6'd55,6'd56,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd59,6'd60,6'd81: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd59,6'd60,6'd61,6'd62,6'd63,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd58,6'd59,6'd60,6'd61,6'd81,6'd82: Enemy_img = 4'd6;
//6'd54,6'd55,6'd84,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd57,6'd58,6'd59,6'd83: Enemy_img = 4'd6;
//6'd51,6'd52,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd57: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd6;
//6'd52,6'd53,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd14;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd14;
//6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72: Enemy_img = 4'd6;
//6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71: Enemy_img = 4'd6;
//6'd72,6'd73: Enemy_img = 4'd7;
//6'd75,6'd76,6'd77,6'd79: Enemy_img = 4'd14;
//6'd78,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71: Enemy_img = 4'd6;
//6'd72,6'd73: Enemy_img = 4'd7;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd82,6'd83,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd6;
//6'd71,6'd72: Enemy_img = 4'd7;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd92,6'd93: Enemy_img = 4'd14;
//6'd81,6'd83,6'd84,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd43,6'd74,6'd75,6'd76,6'd78,6'd80,6'd81,6'd82,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd77,6'd79,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd6;
//6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd93,6'd94: Enemy_img = 4'd13;
//6'd44,6'd75,6'd81,6'd82,6'd83,6'd84,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd49,6'd51,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd6;
//6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd91,6'd92: Enemy_img = 4'd13;
//6'd43,6'd44,6'd73,6'd74,6'd83,6'd84,6'd93,6'd94: Enemy_img = 4'd14;
//6'd45,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd77,6'd78: Enemy_img = 4'd6;
//6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd73,6'd74,6'd86,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd47,6'd75,6'd76,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd78: Enemy_img = 4'd7;
//6'd46,6'd72,6'd73,6'd74,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd44,6'd45,6'd47,6'd75,6'd83,6'd85,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd80: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd44,6'd47,6'd48,6'd83,6'd84,6'd85,6'd89,6'd90: Enemy_img = 4'd14;
//6'd45,6'd46,6'd49,6'd50,6'd73,6'd74,6'd75,6'd82,6'd86,6'd87,6'd88,6'd91,6'd93,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd59,6'd79,6'd80: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd44,6'd45,6'd48,6'd49,6'd73,6'd85,6'd86,6'd87,6'd89,6'd94: Enemy_img = 4'd14;
//6'd46,6'd47,6'd50,6'd72,6'd74,6'd82,6'd83,6'd84,6'd88,6'd90,6'd92,6'd93,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd79,6'd80: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd81: Enemy_img = 4'd7;
//6'd48,6'd49,6'd50,6'd70,6'd71,6'd72,6'd87,6'd88,6'd91,6'd92,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd73,6'd74,6'd75,6'd76,6'd84,6'd85,6'd86,6'd89,6'd90,6'd93,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd78,6'd79: Enemy_img = 4'd6;
//6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd44,6'd46,6'd47,6'd49,6'd71,6'd72,6'd73,6'd74,6'd87,6'd88,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd99,6'd100: Enemy_img = 4'd14;
//6'd43,6'd45,6'd48,6'd50,6'd51,6'd52,6'd53,6'd75,6'd76,6'd77,6'd86,6'd89,6'd98,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd79: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd44,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd107: Enemy_img = 4'd14;
//6'd45,6'd48,6'd49,6'd54,6'd55,6'd56,6'd76,6'd85,6'd106,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd78: Enemy_img = 4'd6;
//6'd62,6'd63,6'd64,6'd65,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd43,6'd44,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//6'd45,6'd47,6'd56,6'd57,6'd58,6'd76,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd42,6'd64,6'd65,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd44,6'd45,6'd52,6'd54,6'd57,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd87,6'd89,6'd90,6'd91,6'd92,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd66,6'd75,6'd84,6'd85,6'd86,6'd88,6'd105,6'd106,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd80,6'd81,6'd82,6'd95: Enemy_img = 4'd6;
//6'd42,6'd94: Enemy_img = 4'd7;
//6'd43,6'd44,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd86,6'd90,6'd91,6'd92,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd45,6'd50,6'd55,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd74,6'd75,6'd76,6'd77,6'd84,6'd85,6'd87,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd81,6'd82,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd41,6'd93,6'd94: Enemy_img = 4'd7;
//6'd43,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd56,6'd58,6'd59,6'd61,6'd70,6'd71,6'd72,6'd74,6'd75,6'd89,6'd90,6'd91,6'd98,6'd99: Enemy_img = 4'd14;
//6'd44,6'd50,6'd54,6'd64,6'd65,6'd66,6'd68,6'd69,6'd73,6'd76,6'd77,6'd78,6'd79,6'd85,6'd86,6'd87,6'd100,6'd101,6'd102,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd82,6'd83,6'd95: Enemy_img = 4'd6;
//6'd41,6'd42,6'd93,6'd94,6'd96: Enemy_img = 4'd7;
//6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd61,6'd64,6'd76,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd43,6'd44,6'd46,6'd50,6'd55,6'd56,6'd57,6'd60,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd85,6'd86,6'd98,6'd99,6'd100,6'd101,6'd103,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd82,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd41,6'd83,6'd96: Enemy_img = 4'd7;
//6'd45,6'd47,6'd51,6'd52,6'd53,6'd56,6'd58,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd89: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49,6'd50,6'd54,6'd55,6'd57,6'd59,6'd60,6'd63,6'd68,6'd69,6'd70,6'd79,6'd86,6'd87,6'd88,6'd99,6'd100,6'd102,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd83,6'd84,6'd85,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd40,6'd41,6'd86,6'd92: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd59,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd47,6'd48,6'd53,6'd58,6'd60,6'd62,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd84,6'd85,6'd86,6'd89,6'd90,6'd92,6'd97: Enemy_img = 4'd6;
//6'd40,6'd41,6'd82,6'd83,6'd87,6'd88,6'd91,6'd94,6'd95,6'd96: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd68,6'd69,6'd71,6'd73,6'd75: Enemy_img = 4'd14;
//6'd47,6'd54,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd70,6'd72,6'd74,6'd76,6'd77,6'd78,6'd79,6'd98,6'd99,6'd100,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd39,6'd40,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd95,6'd96: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd49,6'd50,6'd51,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd71,6'd72,6'd74: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd52,6'd53,6'd62,6'd67,6'd68,6'd69,6'd70,6'd73,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100,6'd101,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd42,6'd43,6'd47,6'd52,6'd53,6'd54,6'd55,6'd57,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd62,6'd70,6'd71,6'd72,6'd91,6'd92,6'd95,6'd96,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd76,6'd77,6'd86,6'd87: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88: Enemy_img = 4'd7;
//6'd42,6'd43,6'd45,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72: Enemy_img = 4'd14;
//6'd21,6'd44,6'd48,6'd49,6'd70,6'd73,6'd74,6'd75,6'd91,6'd94,6'd95,6'd96,6'd97,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd76,6'd77,6'd86,6'd87: Enemy_img = 4'd6;
//6'd37,6'd38,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd64,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd22,6'd23,6'd40,6'd45,6'd49,6'd65,6'd66,6'd67,6'd71,6'd72,6'd93,6'd94,6'd95,6'd96,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd28,6'd30,6'd31,6'd32,6'd33,6'd74,6'd75,6'd86: Enemy_img = 4'd6;
//6'd27,6'd29,6'd34,6'd35,6'd36,6'd37,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd7;
//6'd22,6'd39,6'd40,6'd41,6'd43,6'd44,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd66,6'd67: Enemy_img = 4'd14;
//6'd21,6'd23,6'd42,6'd45,6'd49,6'd64,6'd65,6'd68,6'd69,6'd70,6'd95,6'd97,6'd99,6'd100,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd74,6'd75,6'd76,6'd85,6'd86: Enemy_img = 4'd6;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87: Enemy_img = 4'd7;
//6'd23,6'd24,6'd39,6'd40,6'd41,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd102,6'd103: Enemy_img = 4'd14;
//6'd22,6'd25,6'd42,6'd43,6'd44,6'd45,6'd50,6'd91,6'd92,6'd97,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd86,6'd87: Enemy_img = 4'd6;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd80,6'd81: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd102,6'd103: Enemy_img = 4'd14;
//6'd21,6'd25,6'd46,6'd91,6'd92,6'd93,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73,6'd75,6'd76,6'd78,6'd86,6'd87: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd67,6'd68,6'd69,6'd70,6'd74: Enemy_img = 4'd7;
//6'd103,6'd104: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd102: Enemy_img = 4'd14;
//6'd21,6'd27,6'd37,6'd45,6'd46,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73,6'd87,6'd88: Enemy_img = 4'd6;
//6'd31,6'd68,6'd69,6'd70: Enemy_img = 4'd7;
//6'd102: Enemy_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd39,6'd40,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd103,6'd104: Enemy_img = 4'd14;
//6'd28,6'd35,6'd36,6'd37,6'd38,6'd44,6'd94,6'd95,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60: Enemy_img = 4'd2;
//6'd70,6'd71,6'd87: Enemy_img = 4'd6;
//6'd69,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd42,6'd43,6'd45,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd21,6'd31,6'd37,6'd38,6'd67,6'd77,6'd80,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd2;
//6'd86,6'd87: Enemy_img = 4'd6;
//6'd68,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd63,6'd101,6'd102: Enemy_img = 4'd14;
//6'd21,6'd22,6'd39,6'd64,6'd65,6'd66,6'd75,6'd76,6'd78,6'd79,6'd95,6'd96,6'd97,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd59: Enemy_img = 4'd2;
//6'd86,6'd87: Enemy_img = 4'd6;
//6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd52,6'd53,6'd57,6'd58,6'd61,6'd64,6'd65: Enemy_img = 4'd14;
//6'd62,6'd63,6'd66,6'd70,6'd72,6'd73,6'd74,6'd77,6'd78,6'd83,6'd94,6'd95,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd59: Enemy_img = 4'd2;
//6'd85,6'd86: Enemy_img = 4'd6;
//6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd49: Enemy_img = 4'd9;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd57,6'd62,6'd63: Enemy_img = 4'd14;
//6'd21,6'd61,6'd64,6'd65,6'd66,6'd68,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd96,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd61,6'd62: Enemy_img = 4'd2;
//6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd90: Enemy_img = 4'd7;
//6'd49: Enemy_img = 4'd9;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd56,6'd65: Enemy_img = 4'd14;
//6'd22,6'd57,6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd81,6'd82,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55: Enemy_img = 4'd2;
//6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd48,6'd49: Enemy_img = 4'd9;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd51,6'd52,6'd59,6'd60,6'd64: Enemy_img = 4'd14;
//6'd22,6'd58,6'd65,6'd67,6'd68,6'd69,6'd73,6'd75,6'd76,6'd81,6'd82,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57: Enemy_img = 4'd2;
//6'd92,6'd93: Enemy_img = 4'd6;
//6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd48,6'd49,6'd50: Enemy_img = 4'd10;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd59,6'd60,6'd61,6'd64,6'd65: Enemy_img = 4'd14;
//6'd21,6'd53,6'd62,6'd63,6'd66,6'd69,6'd70,6'd71,6'd75,6'd76,6'd80,6'd83,6'd84,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92: Enemy_img = 4'd6;
//6'd89,6'd90: Enemy_img = 4'd7;
//6'd50: Enemy_img = 4'd9;
//6'd49: Enemy_img = 4'd10;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd53,6'd54,6'd62,6'd64: Enemy_img = 4'd14;
//6'd22,6'd55,6'd60,6'd61,6'd63,6'd65,6'd69,6'd70,6'd73,6'd74,6'd79,6'd80,6'd82,6'd83,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92: Enemy_img = 4'd6;
//6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd50: Enemy_img = 4'd9;
//6'd49: Enemy_img = 4'd10;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55,6'd57,6'd60,6'd62: Enemy_img = 4'd14;
//6'd22,6'd47,6'd56,6'd58,6'd59,6'd61,6'd63,6'd64,6'd65,6'd66,6'd68,6'd71,6'd72,6'd73,6'd74,6'd79,6'd80,6'd81,6'd84,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd91: Enemy_img = 4'd6;
//6'd50: Enemy_img = 4'd9;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd41,6'd42,6'd43,6'd44,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65: Enemy_img = 4'd14;
//6'd22,6'd45,6'd46,6'd47,6'd48,6'd51,6'd56,6'd57,6'd62,6'd63,6'd68,6'd72,6'd73,6'd74,6'd75,6'd79,6'd80,6'd83,6'd84,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd6;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd41,6'd45,6'd46,6'd47,6'd48,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd64: Enemy_img = 4'd14;
//6'd22,6'd42,6'd43,6'd44,6'd51,6'd52,6'd57,6'd58,6'd63,6'd65,6'd68,6'd69,6'd70,6'd73,6'd74,6'd78,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd40: Enemy_img = 4'd6;
//6'd32,6'd35,6'd36,6'd37,6'd38,6'd39: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd55,6'd62,6'd65: Enemy_img = 4'd14;
//6'd42,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd61,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd80,6'd83,6'd85,6'd86,6'd87,6'd90,6'd94,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd40: Enemy_img = 4'd6;
//6'd30,6'd31,6'd35,6'd36,6'd37,6'd38,6'd39,6'd77,6'd79,6'd82,6'd85: Enemy_img = 4'd7;
//6'd23,6'd24,6'd25,6'd26,6'd43,6'd44: Enemy_img = 4'd14;
//6'd22,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd88,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd32,6'd33,6'd38,6'd39: Enemy_img = 4'd6;
//6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd22,6'd23,6'd24,6'd46,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd21,6'd44,6'd45,6'd47,6'd59,6'd61,6'd65,6'd68,6'd72,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd39,6'd40: Enemy_img = 4'd6;
//6'd34,6'd37,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd45,6'd46,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd20,6'd21,6'd41,6'd44,6'd47,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd69,6'd70,6'd92,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd6;
//6'd25,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd47,6'd49: Enemy_img = 4'd14;
//6'd41,6'd46,6'd48,6'd50,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd35,6'd83,6'd85: Enemy_img = 4'd6;
//6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93: Enemy_img = 4'd6;
//6'd26,6'd27,6'd31,6'd32,6'd75,6'd76,6'd77,6'd78,6'd79,6'd92: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd48,6'd49,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd95,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd26,6'd30,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd33,6'd34,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd51,6'd52,6'd54,6'd55,6'd56,6'd60,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd71,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd26,6'd27,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd93,6'd95: Enemy_img = 4'd6;
//6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd51,6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd66,6'd67,6'd70,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd66,6'd69,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd41,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd68,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd25,6'd26,6'd27,6'd28,6'd32,6'd33,6'd37,6'd38,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd72,6'd73: Enemy_img = 4'd7;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd41,6'd44,6'd47,6'd52,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd72,6'd73: Enemy_img = 4'd7;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd60,6'd62,6'd66,6'd67,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd28,6'd29,6'd30,6'd31,6'd36,6'd37,6'd38,6'd39,6'd40,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd51,6'd53,6'd54,6'd72,6'd73,6'd74: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd52,6'd55,6'd56,6'd57: Enemy_img = 4'd7;
//6'd32,6'd33,6'd34,6'd36,6'd37,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd72,6'd73: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd57,6'd58: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd72,6'd73: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd60: Enemy_img = 4'd7;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd56,6'd57,6'd58,6'd59,6'd60,6'd71: Enemy_img = 4'd6;
//6'd42,6'd43: Enemy_img = 4'd7;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd58,6'd59,6'd60,6'd61,6'd62,6'd71: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43: Enemy_img = 4'd7;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd61,6'd62,6'd63,6'd71: Enemy_img = 4'd6;
//6'd41,6'd42: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd64,6'd65: Enemy_img = 4'd6;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd6;
//6'd75: Enemy_img = 4'd7;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd6;
//6'd75: Enemy_img = 4'd7;
//6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73: Enemy_img = 4'd6;
//6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd78,6'd79,6'd80,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd79,6'd81,6'd82,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd6;
//6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd71,6'd72,6'd93,6'd94: Enemy_img = 4'd6;
//6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd92,6'd93: Enemy_img = 4'd6;
//6'd72,6'd73,6'd74,6'd75,6'd76,6'd94: Enemy_img = 4'd7;
//6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd57,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd94,6'd95: Enemy_img = 4'd7;
//6'd48,6'd80,6'd82,6'd84,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd92,6'd97: Enemy_img = 4'd6;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd7;
//6'd49,6'd50,6'd76,6'd78,6'd84,6'd86,6'd87,6'd88,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd91,6'd92,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd89,6'd90,6'd93,6'd94: Enemy_img = 4'd7;
//6'd99,6'd100: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd75,6'd76,6'd77,6'd79,6'd80,6'd82,6'd83,6'd86,6'd87,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd98,6'd99: Enemy_img = 4'd14;
//6'd50,6'd52,6'd54,6'd55,6'd57,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95: Enemy_img = 4'd6;
//6'd63,6'd64,6'd65,6'd66,6'd87,6'd88,6'd94: Enemy_img = 4'd7;
//6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd51,6'd52,6'd54,6'd57,6'd58,6'd60,6'd66,6'd68,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd88,6'd92,6'd93: Enemy_img = 4'd7;
//6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd78,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd84,6'd85,6'd90: Enemy_img = 4'd6;
//6'd86,6'd87,6'd88,6'd89,6'd91,6'd92: Enemy_img = 4'd7;
//6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd62,6'd65,6'd66,6'd69,6'd70,6'd71,6'd80,6'd81,6'd82,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd83,6'd84,6'd89,6'd90: Enemy_img = 4'd6;
//6'd85,6'd86,6'd87,6'd88,6'd91: Enemy_img = 4'd7;
//6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd68,6'd69,6'd70,6'd71,6'd73,6'd81,6'd82,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd84,6'd89,6'd90: Enemy_img = 4'd6;
//6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd74,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd83,6'd84,6'd88,6'd89: Enemy_img = 4'd6;
//6'd49,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd74,6'd76,6'd78,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd52,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd73,6'd75,6'd77,6'd79,6'd81,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd49: Enemy_img = 4'd7;
//6'd74,6'd75,6'd77,6'd78,6'd80,6'd90,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd53,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd76,6'd79,6'd81,6'd82,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd85,6'd87: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50: Enemy_img = 4'd7;
//6'd74,6'd75,6'd79,6'd80,6'd81,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd53,6'd54,6'd58,6'd59,6'd60,6'd62,6'd63,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48: Enemy_img = 4'd6;
//6'd49,6'd50: Enemy_img = 4'd7;
//6'd74,6'd77,6'd78,6'd79,6'd80,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd53,6'd56,6'd57,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd73,6'd75,6'd76,6'd81,6'd82,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47: Enemy_img = 4'd6;
//6'd48,6'd49: Enemy_img = 4'd7;
//6'd76,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd14;
//6'd53,6'd54,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd73,6'd74,6'd75,6'd80,6'd81,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50: Enemy_img = 4'd7;
//6'd75,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd53,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd74,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50: Enemy_img = 4'd7;
//6'd75: Enemy_img = 4'd9;
//6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd70,6'd71,6'd74,6'd78,6'd79,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd7;
//6'd76: Enemy_img = 4'd9;
//6'd70,6'd71,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd69,6'd73,6'd75,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd7;
//6'd76: Enemy_img = 4'd9;
//6'd77: Enemy_img = 4'd10;
//6'd70,6'd71,6'd72,6'd73,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd102,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd66,6'd68,6'd69,6'd98,6'd101,6'd103,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd77,6'd78: Enemy_img = 4'd10;
//6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92,6'd94,6'd106,6'd107: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd93,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd7;
//6'd78,6'd79: Enemy_img = 4'd9;
//6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd73,6'd75,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd90: Enemy_img = 4'd14;
//6'd55,6'd57,6'd58,6'd62,6'd68,6'd69,6'd70,6'd71,6'd74,6'd89,6'd91,6'd92,6'd93,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd101,6'd102,6'd103: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd79: Enemy_img = 4'd9;
//6'd62,6'd64,6'd66,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd14;
//6'd53,6'd54,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd65,6'd67,6'd68,6'd71,6'd74,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd2;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd78: Enemy_img = 4'd9;
//6'd62,6'd63,6'd75,6'd76,6'd77,6'd81,6'd82,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd2;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd94,6'd95,6'd96: Enemy_img = 4'd7;
//6'd62,6'd65,6'd67,6'd68,6'd75,6'd76,6'd77,6'd80,6'd82,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd55,6'd57,6'd58,6'd61,6'd63,6'd64,6'd66,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd2;
//6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd93,6'd94,6'd95: Enemy_img = 4'd7;
//6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd59,6'd62,6'd65,6'd70,6'd71,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd69,6'd73: Enemy_img = 4'd2;
//6'd30,6'd32,6'd33,6'd34,6'd36,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd63,6'd64,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd26,6'd28,6'd53,6'd54,6'd55,6'd56,6'd62,6'd83,6'd84,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70: Enemy_img = 4'd2;
//6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd64,6'd71,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd85,6'd89,6'd90: Enemy_img = 4'd14;
//6'd27,6'd30,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd62,6'd63,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd36,6'd38,6'd39,6'd41,6'd42,6'd92,6'd93: Enemy_img = 4'd7;
//6'd63,6'd66,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88: Enemy_img = 4'd14;
//6'd28,6'd31,6'd32,6'd33,6'd44,6'd48,6'd49,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd67,6'd68,6'd85,6'd86,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd92,6'd93: Enemy_img = 4'd7;
//6'd65,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd54,6'd57,6'd60,6'd61,6'd63,6'd64,6'd66,6'd67,6'd80,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70: Enemy_img = 4'd2;
//6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd91,6'd92: Enemy_img = 4'd7;
//6'd64,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd53,6'd55,6'd56,6'd58,6'd59,6'd61,6'd65,6'd66,6'd81,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd91,6'd92: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd35,6'd38,6'd42,6'd44,6'd45,6'd48,6'd49,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd64,6'd65,6'd82,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd62,6'd91,6'd92: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd31,6'd46,6'd47,6'd49,6'd53,6'd54,6'd55,6'd57,6'd58,6'd63,6'd83,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd93,6'd94: Enemy_img = 4'd6;
//6'd39,6'd61,6'd62,6'd91,6'd92: Enemy_img = 4'd7;
//6'd64,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd32,6'd34,6'd45,6'd46,6'd48,6'd53,6'd54,6'd56,6'd57,6'd82,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd60,6'd93,6'd94: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd61,6'd62,6'd63,6'd64,6'd92: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd45,6'd48,6'd49,6'd53,6'd55,6'd56,6'd81,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd59,6'd93,6'd94: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd60,6'd61,6'd62,6'd63,6'd92: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd34,6'd48,6'd52,6'd55,6'd80,6'd86,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd41,6'd42,6'd45,6'd59,6'd60,6'd62,6'd93,6'd94: Enemy_img = 4'd6;
//6'd40,6'd58,6'd61: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd70,6'd72,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd88,6'd90: Enemy_img = 4'd14;
//6'd32,6'd48,6'd52,6'd53,6'd68,6'd79,6'd85,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd58,6'd59,6'd60,6'd61,6'd93,6'd94: Enemy_img = 4'd6;
//6'd57,6'd92: Enemy_img = 4'd7;
//6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd76,6'd78,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd91: Enemy_img = 4'd14;
//6'd33,6'd34,6'd51,6'd64,6'd67,6'd79,6'd80,6'd84,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd54,6'd56,6'd57,6'd58,6'd59,6'd93,6'd94: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd60: Enemy_img = 4'd7;
//6'd64,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd85,6'd86,6'd87,6'd90,6'd91: Enemy_img = 4'd14;
//6'd33,6'd34,6'd63,6'd65,6'd66,6'd71,6'd80,6'd83,6'd84,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd59: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd74,6'd75,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd33,6'd34,6'd62,6'd73,6'd76,6'd79,6'd84,6'd85,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd53,6'd54,6'd57,6'd58,6'd94: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd52,6'd55,6'd56: Enemy_img = 4'd7;
//6'd62,6'd64,6'd65,6'd67,6'd68,6'd70,6'd73,6'd76,6'd79,6'd81,6'd82,6'd91: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd61,6'd63,6'd66,6'd69,6'd71,6'd72,6'd74,6'd75,6'd77,6'd78,6'd80,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd57,6'd94: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd46,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd7;
//6'd61,6'd62,6'd64,6'd70,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd35,6'd37,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd74,6'd82,6'd84,6'd86,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd56,6'd57,6'd58,6'd94,6'd95: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd7;
//6'd60,6'd61,6'd66,6'd69,6'd70,6'd73,6'd74,6'd76,6'd81,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90: Enemy_img = 4'd14;
//6'd36,6'd37,6'd59,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd72,6'd75,6'd80,6'd82,6'd87,6'd88,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd56,6'd57: Enemy_img = 4'd6;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd7;
//6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd92,6'd93: Enemy_img = 4'd14;
//6'd29,6'd31,6'd34,6'd35,6'd36,6'd59,6'd61,6'd62,6'd64,6'd76,6'd78,6'd86,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd7;
//6'd31,6'd32,6'd60,6'd61,6'd86,6'd87,6'd88,6'd92,6'd93: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd7;
//6'd30,6'd31,6'd59,6'd87,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd69,6'd70,6'd73,6'd75,6'd76,6'd79,6'd80,6'd82,6'd83,6'd85,6'd86,6'd88,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd28,6'd40,6'd56,6'd57,6'd58,6'd59,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd86: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd31,6'd32: Enemy_img = 4'd13;
//6'd29,6'd30,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd94: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd59,6'd61,6'd63,6'd70,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd50,6'd51,6'd53,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd91: Enemy_img = 4'd6;
//6'd48,6'd49,6'd52,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd7;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd95: Enemy_img = 4'd14;
//6'd34,6'd37,6'd39,6'd40,6'd41,6'd44,6'd55,6'd57,6'd58,6'd59,6'd63,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd31,6'd32,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd35,6'd39,6'd40,6'd41,6'd43,6'd44,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd54,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd45,6'd47,6'd50,6'd51,6'd53,6'd55,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd32,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd43,6'd57,6'd58,6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd46,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76: Enemy_img = 4'd7;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd48,6'd49,6'd50,6'd51,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd55,6'd56,6'd58,6'd59,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd57,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd47,6'd48,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd50,6'd51,6'd52,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd41,6'd42,6'd43,6'd59,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd40,6'd44,6'd55,6'd56,6'd57,6'd58,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd46,6'd47,6'd48,6'd51,6'd64,6'd66,6'd67: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd50,6'd52,6'd53,6'd61,6'd62,6'd63,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd59,6'd60,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd44,6'd55,6'd56,6'd57,6'd58,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd65,6'd66: Enemy_img = 4'd14;
//6'd36,6'd37,6'd50,6'd52,6'd53,6'd61,6'd62,6'd63,6'd64,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd42,6'd43,6'd59,6'd60,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd41,6'd44,6'd55,6'd56,6'd57,6'd58,6'd61,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd46,6'd47,6'd48,6'd67: Enemy_img = 4'd14;
//6'd34,6'd50,6'd51,6'd52,6'd53,6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd59,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd43,6'd44,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd46,6'd47,6'd48,6'd52,6'd66: Enemy_img = 4'd14;
//6'd33,6'd34,6'd38,6'd39,6'd50,6'd51,6'd53,6'd54,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd43,6'd59,6'd60,6'd72,6'd73,6'd74: Enemy_img = 4'd6;
//6'd44,6'd61,6'd62,6'd63,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd40,6'd46,6'd47,6'd48,6'd51,6'd52,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd50,6'd53,6'd55,6'd56,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd63,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd6;
//6'd62,6'd68,6'd69,6'd70: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd43,6'd44,6'd46,6'd47,6'd48,6'd51,6'd52,6'd66,6'd67: Enemy_img = 4'd14;
//6'd34,6'd37,6'd38,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd62,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd69,6'd70: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd55,6'd56: Enemy_img = 4'd14;
//6'd33,6'd36,6'd37,6'd50,6'd51,6'd54,6'd57,6'd58,6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd6;
//6'd68,6'd69: Enemy_img = 4'd7;
//6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd56,6'd66,6'd67: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd37,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd6;
//6'd69,6'd70: Enemy_img = 4'd7;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd51,6'd54,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd33,6'd34,6'd47,6'd50,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd6;
//6'd69: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd52,6'd53,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd33,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd56,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd32,6'd38,6'd39,6'd41,6'd42,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71: Enemy_img = 4'd6;
//6'd33,6'd49,6'd52,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd32,6'd34,6'd36,6'd37,6'd46,6'd47,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50: Enemy_img = 4'd13;
//6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd62,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd31,6'd32,6'd59,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71: Enemy_img = 4'd6;
//6'd49: Enemy_img = 4'd13;
//6'd48,6'd50,6'd51,6'd52,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd67: Enemy_img = 4'd14;
//6'd52,6'd53,6'd64,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd68,6'd70: Enemy_img = 4'd14;
//6'd51,6'd52,6'd67,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd14;
//6'd51,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70: Enemy_img = 4'd14;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd60,6'd61,6'd63,6'd64,6'd66,6'd69,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd77: Enemy_img = 4'd6;
//6'd78: Enemy_img = 4'd7;
//6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd74,6'd75,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd77,6'd78,6'd82: Enemy_img = 4'd6;
//6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd84: Enemy_img = 4'd14;
//6'd61,6'd62,6'd63,6'd64,6'd69,6'd70,6'd71,6'd74,6'd75,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd76,6'd77,6'd78,6'd81,6'd82: Enemy_img = 4'd6;
//6'd58,6'd59,6'd79,6'd80: Enemy_img = 4'd7;
//6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd6;
//6'd59,6'd60,6'd76,6'd79: Enemy_img = 4'd7;
//6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd63,6'd65,6'd66,6'd67,6'd71,6'd73,6'd74,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd61,6'd76: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd65,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd75,6'd76,6'd81: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd77,6'd78: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62,6'd75,6'd76,6'd79,6'd80: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd64,6'd65,6'd66,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd74,6'd79,6'd80: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd69,6'd71,6'd72,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd79: Enemy_img = 4'd7;
//6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd66,6'd71,6'd72,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd74,6'd75,6'd78: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd61,6'd76,6'd77,6'd79: Enemy_img = 4'd7;
//6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd63,6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd73,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd73,6'd77,6'd78: Enemy_img = 4'd6;
//6'd58,6'd59,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd61,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd72,6'd73,6'd78: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd72,6'd73,6'd76,6'd77: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd74,6'd75: Enemy_img = 4'd7;
//6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd69,6'd70,6'd71,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd73,6'd76,6'd77: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd74,6'd75: Enemy_img = 4'd7;
//6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd94,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd74,6'd75,6'd77: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd7;
//6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd90: Enemy_img = 4'd14;
//6'd57,6'd59,6'd60,6'd61,6'd89,6'd91,6'd92,6'd93,6'd95,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd96: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd91,6'd93,6'd94: Enemy_img = 4'd7;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd57,6'd59,6'd60,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd45,6'd95: Enemy_img = 4'd6;
//6'd47,6'd48,6'd50,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd63,6'd65,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95: Enemy_img = 4'd6;
//6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd64,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd36,6'd38,6'd44,6'd46,6'd48,6'd49,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd63,6'd65,6'd66,6'd67,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92,6'd93: Enemy_img = 4'd6;
//6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd65,6'd66,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd55,6'd56,6'd60,6'd61,6'd62,6'd64,6'd67,6'd68,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92,6'd93: Enemy_img = 4'd6;
//6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd65,6'd66,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd39,6'd40,6'd43,6'd44,6'd47,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd61,6'd67,6'd71,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd65,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd83: Enemy_img = 4'd14;
//6'd39,6'd44,6'd46,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd61,6'd62,6'd66,6'd71,6'd82,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd88,6'd89: Enemy_img = 4'd7;
//6'd67,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd45,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd61,6'd62,6'd65,6'd66,6'd70,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd87,6'd88: Enemy_img = 4'd7;
//6'd68,6'd69: Enemy_img = 4'd9;
//6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd61,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd87,6'd88: Enemy_img = 4'd7;
//6'd68: Enemy_img = 4'd9;
//6'd69,6'd70,6'd71: Enemy_img = 4'd10;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd50,6'd54,6'd56,6'd57,6'd58,6'd64,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd90,6'd91: Enemy_img = 4'd6;
//6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd69,6'd71,6'd72: Enemy_img = 4'd9;
//6'd70: Enemy_img = 4'd10;
//6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd43,6'd44,6'd46,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd87,6'd88: Enemy_img = 4'd7;
//6'd72,6'd73: Enemy_img = 4'd9;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd74,6'd75,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd44,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd90,6'd91: Enemy_img = 4'd6;
//6'd41,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd73: Enemy_img = 4'd9;
//6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd75,6'd77,6'd78,6'd80,6'd81,6'd85: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd68,6'd79,6'd82,6'd83,6'd84,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd41,6'd42,6'd87,6'd88: Enemy_img = 4'd7;
//6'd62,6'd66,6'd67,6'd69,6'd70,6'd71,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd83,6'd85: Enemy_img = 4'd14;
//6'd45,6'd46,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd63,6'd64,6'd65,6'd79,6'd82,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd2;
//6'd39,6'd40,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd87,6'd88: Enemy_img = 4'd7;
//6'd61,6'd62,6'd64,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd63,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd68: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd90,6'd91: Enemy_img = 4'd6;
//6'd42,6'd43,6'd88,6'd89: Enemy_img = 4'd7;
//6'd59,6'd60,6'd61,6'd62,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd46,6'd50,6'd53,6'd57,6'd58,6'd63,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd88,6'd89: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd61,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd56,6'd57,6'd62,6'd67,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd91,6'd92: Enemy_img = 4'd6;
//6'd42,6'd43,6'd89,6'd90: Enemy_img = 4'd7;
//6'd56,6'd63,6'd64,6'd67,6'd71,6'd72,6'd73,6'd74,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86: Enemy_img = 4'd14;
//6'd47,6'd50,6'd51,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd77,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd90: Enemy_img = 4'd7;
//6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd81,6'd82,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd53,6'd56,6'd59,6'd78,6'd79,6'd80,6'd83,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd42,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45: Enemy_img = 4'd7;
//6'd58,6'd62,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd49,6'd50,6'd52,6'd53,6'd57,6'd59,6'd60,6'd61,6'd80,6'd81,6'd82,6'd83,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd92,6'd93: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd91: Enemy_img = 4'd7;
//6'd59,6'd60,6'd61,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd57,6'd58,6'd80,6'd83,6'd84,6'd85,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd93,6'd94: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd7;
//6'd59,6'd60,6'd61,6'd63,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd89,6'd90: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd64,6'd65,6'd80,6'd84,6'd85,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd2;
//6'd38,6'd39,6'd40,6'd93,6'd94: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd61,6'd63,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd51,6'd59,6'd60,6'd62,6'd64,6'd79,6'd84,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd94: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd63,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd58,6'd60,6'd61,6'd62,6'd64,6'd79,6'd83,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd95: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd80,6'd81,6'd82,6'd85,6'd89: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd54,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd78,6'd79,6'd83,6'd84,6'd88,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd95: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd55,6'd58,6'd59,6'd60,6'd62,6'd63,6'd79,6'd80,6'd85,6'd87,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd71,6'd76,6'd78,6'd79,6'd81,6'd82,6'd83,6'd86,6'd87,6'd90,6'd91,6'd93,6'd94: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd57,6'd62,6'd80,6'd85,6'd88,6'd89,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd61: Enemy_img = 4'd7;
//6'd63,6'd67,6'd68,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82,6'd86,6'd87,6'd96: Enemy_img = 4'd14;
//6'd47,6'd54,6'd57,6'd58,6'd59,6'd79,6'd80,6'd81,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd61,6'd62,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd80,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd52,6'd55,6'd56,6'd57,6'd77,6'd78,6'd79,6'd81,6'd83,6'd88,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd60: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd61,6'd62,6'd63: Enemy_img = 4'd7;
//6'd66,6'd67,6'd69,6'd70,6'd73,6'd77,6'd78,6'd80,6'd83,6'd84,6'd85,6'd86,6'd89,6'd92,6'd94,6'd97,6'd98: Enemy_img = 4'd14;
//6'd47,6'd48,6'd52,6'd53,6'd54,6'd57,6'd68,6'd71,6'd72,6'd74,6'd75,6'd76,6'd79,6'd82,6'd87,6'd88,6'd90,6'd91,6'd93,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd60,6'd63: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd61,6'd62: Enemy_img = 4'd7;
//6'd65,6'd66,6'd68,6'd69,6'd70,6'd73,6'd75,6'd77,6'd78,6'd82,6'd84: Enemy_img = 4'd14;
//6'd43,6'd45,6'd47,6'd48,6'd49,6'd52,6'd53,6'd54,6'd56,6'd57,6'd67,6'd74,6'd76,6'd80,6'd81,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd59,6'd60,6'd61,6'd62,6'd63,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd88: Enemy_img = 4'd7;
//6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd78,6'd81: Enemy_img = 4'd14;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd53,6'd54,6'd56,6'd65,6'd66,6'd67,6'd73,6'd76,6'd77,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd60,6'd61,6'd62,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd59,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd75,6'd76: Enemy_img = 4'd14;
//6'd40,6'd42,6'd43,6'd44,6'd45,6'd49,6'd53,6'd54,6'd56,6'd64,6'd71,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd31,6'd60,6'd61,6'd62,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd33,6'd34,6'd36,6'd58,6'd59,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd44,6'd47,6'd49,6'd53,6'd64,6'd68,6'd69,6'd70,6'd75,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd61,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd67,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd30,6'd32,6'd35,6'd36,6'd37,6'd41,6'd46,6'd49,6'd54,6'd55,6'd63,6'd64,6'd65,6'd66,6'd68,6'd70,6'd74,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd64,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38,6'd45,6'd46,6'd49,6'd53,6'd63,6'd65,6'd66,6'd67,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd59,6'd60,6'd61,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd42,6'd58,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd64,6'd66,6'd68,6'd69: Enemy_img = 4'd14;
//6'd28,6'd29,6'd31,6'd32,6'd35,6'd36,6'd50,6'd63,6'd65,6'd67,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd47,6'd56,6'd57,6'd60,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd41,6'd42,6'd58,6'd59,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd63,6'd67: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd62,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd44,6'd46,6'd47,6'd60,6'd61,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd55,6'd56,6'd57,6'd58,6'd59,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd64,6'd65,6'd73: Enemy_img = 4'd14;
//6'd32,6'd33,6'd36,6'd63,6'd66,6'd67,6'd70,6'd71,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd42,6'd43,6'd44,6'd45,6'd47,6'd60,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd41,6'd46,6'd55,6'd56,6'd57,6'd58,6'd59,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd64,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd32,6'd34,6'd35,6'd36,6'd62,6'd63,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd48,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd63,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd62,6'd64,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd48,6'd49,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd34,6'd62,6'd63,6'd64,6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd67,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd61,6'd62,6'd64,6'd65,6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd52,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd37,6'd38,6'd61,6'd64,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd44,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd60,6'd63,6'd64,6'd65,6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd59,6'd66,6'd67,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd70,6'd71,6'd73: Enemy_img = 4'd14;
//6'd38,6'd39,6'd42,6'd62,6'd63,6'd68,6'd69,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd52,6'd54,6'd55,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd73: Enemy_img = 4'd14;
//6'd41,6'd45,6'd47,6'd48,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd58,6'd59,6'd66,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd74: Enemy_img = 4'd14;
//6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd62,6'd67,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd63,6'd64,6'd65,6'd66,6'd71,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd74,6'd75: Enemy_img = 4'd14;
//6'd40,6'd43,6'd44,6'd45,6'd46,6'd50,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd67,6'd68,6'd80,6'd81: Enemy_img = 4'd6;
//6'd54,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd75,6'd76: Enemy_img = 4'd14;
//6'd37,6'd41,6'd42,6'd47,6'd51,6'd57,6'd58,6'd59,6'd60,6'd61,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd68,6'd80,6'd81: Enemy_img = 4'd6;
//6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd37,6'd76: Enemy_img = 4'd14;
//6'd35,6'd36,6'd41,6'd46,6'd47,6'd48,6'd50,6'd56,6'd58,6'd59,6'd60,6'd61,6'd73,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd68,6'd70,6'd71,6'd72,6'd80,6'd81: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66,6'd69,6'd79: Enemy_img = 4'd7;
//6'd37,6'd38,6'd55,6'd56,6'd59,6'd60,6'd75,6'd76: Enemy_img = 4'd14;
//6'd35,6'd36,6'd43,6'd44,6'd47,6'd48,6'd61,6'd62,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd69,6'd70,6'd71,6'd81: Enemy_img = 4'd6;
//6'd64,6'd79,6'd80: Enemy_img = 4'd7;
//6'd39: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd55,6'd56,6'd57,6'd59,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd34,6'd35,6'd42,6'd46,6'd47,6'd48,6'd58,6'd60,6'd61,6'd62,6'd63,6'd67,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd69,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd49,6'd50: Enemy_img = 4'd7;
//6'd38: Enemy_img = 4'd13;
//6'd36,6'd37,6'd39,6'd54,6'd55,6'd56,6'd57,6'd61,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd35,6'd42,6'd43,6'd44,6'd46,6'd59,6'd60,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd81: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd53: Enemy_img = 4'd7;
//6'd38: Enemy_img = 4'd13;
//6'd37,6'd39,6'd40,6'd55,6'd56,6'd57,6'd61,6'd62,6'd65,6'd66,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd59,6'd60,6'd63,6'd64,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd82: Enemy_img = 4'd6;
//6'd53,6'd54: Enemy_img = 4'd7;
//6'd39,6'd40,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd41,6'd43,6'd44,6'd45,6'd46,6'd64,6'd65,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd52: Enemy_img = 4'd6;
//6'd50,6'd51,6'd53,6'd54: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd76,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd52,6'd53: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd73,6'd78,6'd79,6'd82: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd60,6'd63,6'd64,6'd67,6'd72,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd81,6'd82: Enemy_img = 4'd14;
//6'd48,6'd49,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd62,6'd83: Enemy_img = 4'd14;
//6'd44,6'd45,6'd48,6'd49,6'd58,6'd59,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd14;
//6'd44,6'd46,6'd47,6'd48,6'd59,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd64,6'd65: Enemy_img = 4'd14;
//6'd45,6'd48,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd60,6'd61,6'd62,6'd64,6'd65: Enemy_img = 4'd14;
//6'd48,6'd49,6'd54,6'd55,6'd56,6'd58,6'd59,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd45,6'd47,6'd55,6'd59,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd52,6'd53,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd64: Enemy_img = 4'd14;
//6'd45,6'd46,6'd51,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd14;
//6'd46,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd14;
//6'd45,6'd46,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd64: Enemy_img = 4'd6;
//6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd64: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd56,6'd57,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd56,6'd57,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd59,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd56,6'd57,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd59,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd56,6'd57,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd53,6'd54,6'd56,6'd57,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd54,6'd56,6'd57,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd59,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd54,6'd56,6'd57,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd60,6'd61,6'd62,6'd63,6'd82: Enemy_img = 4'd6;
//6'd59,6'd64: Enemy_img = 4'd7;
//6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd54,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd59,6'd60,6'd63,6'd64,6'd82: Enemy_img = 4'd6;
//6'd42,6'd43,6'd61,6'd62,6'd80,6'd81: Enemy_img = 4'd7;
//6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd56,6'd57,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd59,6'd60,6'd63,6'd64,6'd81,6'd82: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd61,6'd62,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd54,6'd56,6'd57,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd59,6'd64,6'd81: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd60,6'd61,6'd62,6'd63,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74: Enemy_img = 4'd14;
//6'd49,6'd56,6'd57,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd59,6'd64,6'd80,6'd81: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd60,6'd61,6'd62,6'd63,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd50,6'd52,6'd53,6'd54,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd59,6'd60,6'd63,6'd64,6'd80,6'd81: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd61,6'd62,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd59,6'd60,6'd63,6'd64,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd61,6'd62,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd60,6'd61,6'd62,6'd63,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd54,6'd56,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd46,6'd77,6'd78: Enemy_img = 4'd7;
//6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75: Enemy_img = 4'd14;
//6'd48,6'd49,6'd59,6'd60,6'd61,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd46,6'd77,6'd78: Enemy_img = 4'd7;
//6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd74,6'd75: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd61,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd58,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd44,6'd45,6'd78,6'd79: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd53,6'd54,6'd58,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd53,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd48,6'd49,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd43,6'd44,6'd79,6'd80: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49,6'd50,6'd53,6'd57,6'd61,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd55,6'd56,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd77: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49,6'd50,6'd51,6'd54,6'd57,6'd60,6'd61,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd56,6'd58,6'd65,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd55,6'd57,6'd71,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd59,6'd60,6'd64: Enemy_img = 4'd9;
//6'd61,6'd62,6'd63: Enemy_img = 4'd10;
//6'd66,6'd67,6'd69,6'd70,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd52,6'd53,6'd56,6'd57,6'd71,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd39,6'd40,6'd83,6'd84: Enemy_img = 4'd7;
//6'd60,6'd61,6'd63,6'd64,6'd65: Enemy_img = 4'd9;
//6'd62: Enemy_img = 4'd10;
//6'd67,6'd69,6'd70,6'd78,6'd79: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd52,6'd53,6'd56,6'd58,6'd59,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd38,6'd85: Enemy_img = 4'd7;
//6'd65: Enemy_img = 4'd9;
//6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd49,6'd50,6'd52,6'd53,6'd56,6'd58,6'd77,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd83,6'd84: Enemy_img = 4'd14;
//6'd39,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd52,6'd53,6'd56,6'd77,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd89,6'd90: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd55,6'd61,6'd77,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd91: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd55,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd2;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd89,6'd90: Enemy_img = 4'd14;
//6'd33,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd75,6'd79,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd63: Enemy_img = 4'd2;
//6'd56,6'd58,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87,6'd89,6'd90,6'd92,6'd93: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd41,6'd49,6'd50,6'd51,6'd52,6'd55,6'd57,6'd75,6'd79,6'd84,6'd88,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd64: Enemy_img = 4'd2;
//6'd55,6'd56,6'd62,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd57,6'd61,6'd75,6'd79,6'd83,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd84,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd57,6'd60,6'd61,6'd75,6'd79,6'd80,6'd81,6'd83,6'd85,6'd86,6'd87,6'd88,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd47,6'd48,6'd49,6'd50,6'd53,6'd57,6'd75,6'd82,6'd85,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd2;
//6'd31,6'd92: Enemy_img = 4'd6;
//6'd53,6'd54,6'd58,6'd59,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd78,6'd79,6'd80,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd52,6'd55,6'd56,6'd57,6'd75,6'd76,6'd77,6'd82,6'd85,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd63: Enemy_img = 4'd2;
//6'd32,6'd33,6'd90,6'd91: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd78,6'd79,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd38,6'd40,6'd41,6'd44,6'd45,6'd47,6'd48,6'd51,6'd52,6'd53,6'd54,6'd55,6'd77,6'd81,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd64: Enemy_img = 4'd2;
//6'd33,6'd34,6'd89,6'd90: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd62,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd82,6'd83: Enemy_img = 4'd14;
//6'd40,6'd41,6'd44,6'd45,6'd50,6'd51,6'd55,6'd56,6'd57,6'd61,6'd77,6'd78,6'd79,6'd81,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd36,6'd87: Enemy_img = 4'd7;
//6'd54,6'd56,6'd57,6'd60,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd76,6'd78,6'd81,6'd82: Enemy_img = 4'd14;
//6'd41,6'd42,6'd45,6'd46,6'd47,6'd52,6'd53,6'd55,6'd61,6'd77,6'd80,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd88,6'd89: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd56,6'd57,6'd58,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd78,6'd81: Enemy_img = 4'd14;
//6'd42,6'd45,6'd46,6'd47,6'd49,6'd54,6'd55,6'd59,6'd61,6'd75,6'd76,6'd77,6'd80,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd58,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd80: Enemy_img = 4'd14;
//6'd43,6'd46,6'd47,6'd49,6'd50,6'd51,6'd56,6'd57,6'd59,6'd61,6'd75,6'd79,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd60,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd76,6'd77: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd58,6'd59,6'd61,6'd73,6'd74,6'd75,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd41,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd62,6'd63,6'd66,6'd67,6'd72,6'd74: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd56,6'd57,6'd60,6'd61,6'd70,6'd71,6'd73,6'd75,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd62,6'd65,6'd66,6'd68,6'd69,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd67,6'd72,6'd73,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd60,6'd63,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd65,6'd66,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd52,6'd54,6'd67,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd60,6'd61,6'd62,6'd63,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd65,6'd66,6'd68,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd54,6'd56,6'd57,6'd58,6'd67,6'd71,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd60,6'd63,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd61,6'd62,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd68,6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd56,6'd57,6'd65,6'd66,6'd67,6'd71,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd60,6'd63,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd61,6'd62,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd72,6'd73: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd65,6'd69,6'd70,6'd71,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd60,6'd61,6'd62,6'd63,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd57,6'd65,6'd69,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd60,6'd61,6'd62,6'd63,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd68,6'd70,6'd71: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd57,6'd65,6'd66,6'd67,6'd69,6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd61,6'd62,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd60,6'd63,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd66,6'd70,6'd75,6'd76: Enemy_img = 4'd14;
//6'd47,6'd48,6'd53,6'd54,6'd55,6'd57,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd61,6'd62,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd60,6'd63,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd66,6'd68,6'd69,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd49,6'd54,6'd55,6'd57,6'd65,6'd67,6'd70,6'd71,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd60,6'd61,6'd62,6'd63,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd66,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd55,6'd65,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd60,6'd61,6'd62,6'd63,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd46,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57,6'd65,6'd69,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd59,6'd60,6'd63,6'd64,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd61,6'd62,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd45,6'd46,6'd51,6'd56,6'd66,6'd68,6'd69,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd59,6'd60,6'd63,6'd64,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd61,6'd62,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd67,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd49,6'd51,6'd52,6'd56,6'd66,6'd68,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd59,6'd64,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd60,6'd61,6'd62,6'd63,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd49,6'd52,6'd66,6'd67,6'd68,6'd70,6'd72,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd86,6'd87: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd41,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd70,6'd74,6'd75,6'd76,6'd78,6'd80: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd49,6'd53,6'd66,6'd67,6'd69,6'd71,6'd72,6'd73,6'd77,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd75,6'd80,6'd81: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd48,6'd66,6'd67,6'd69,6'd70,6'd71,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd51,6'd72,6'd87,6'd88: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd66,6'd68,6'd69,6'd70,6'd74,6'd75,6'd76,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd50,6'd51,6'd52,6'd71,6'd72,6'd73,6'd88,6'd89: Enemy_img = 4'd6;
//6'd36,6'd37,6'd46,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd77,6'd86,6'd87: Enemy_img = 4'd7;
//6'd83: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd66,6'd68,6'd69,6'd75,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd49,6'd50,6'd52,6'd53,6'd70,6'd71,6'd73,6'd74,6'd88,6'd89: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd51,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd72,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd44,6'd48,6'd49,6'd53,6'd54,6'd56,6'd57,6'd58,6'd65,6'd66,6'd67,6'd69,6'd70,6'd74,6'd75,6'd79,6'd90: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd50,6'd51,6'd52,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd68,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd36,6'd37,6'd39,6'd40,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd47,6'd48,6'd54,6'd55,6'd56,6'd58,6'd59,6'd64,6'd65,6'd67,6'd68,6'd69,6'd75,6'd76,6'd78,6'd79: Enemy_img = 4'd6;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd60,6'd61,6'd62,6'd63,6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd77: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd59,6'd60,6'd63,6'd64,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd58,6'd61,6'd62,6'd65,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91: Enemy_img = 4'd14;
//6'd32,6'd36,6'd37,6'd38,6'd39,6'd41,6'd80,6'd81,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd60,6'd63,6'd77: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd59,6'd61,6'd62,6'd64,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd41,6'd42,6'd66,6'd67,6'd68,6'd69,6'd75,6'd79,6'd80,6'd81,6'd85,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd51,6'd60,6'd63,6'd72: Enemy_img = 4'd7;
//6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd38,6'd40,6'd41,6'd42,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd75,6'd76,6'd78,6'd79,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd6;
//6'd62: Enemy_img = 4'd7;
//6'd67,6'd68,6'd75,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd14;
//6'd40,6'd44,6'd54,6'd55,6'd56,6'd64,6'd66,6'd69,6'd70,6'd71,6'd73,6'd74,6'd76,6'd77,6'd78,6'd82,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd64,6'd65,6'd68,6'd70,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd49,6'd53,6'd54,6'd55,6'd58,6'd59,6'd67,6'd69,6'd71,6'd72,6'd73,6'd77,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd6;
//6'd61: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd70,6'd71,6'd73,6'd78,6'd79: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd49,6'd52,6'd53,6'd54,6'd59,6'd68,6'd69,6'd72,6'd74,6'd75,6'd76,6'd77,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd46,6'd49,6'd51,6'd52,6'd53,6'd56,6'd57,6'd59,6'd69,6'd74,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd6;
//6'd62: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd75: Enemy_img = 4'd14;
//6'd48,6'd49,6'd55,6'd56,6'd57,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd60,6'd63: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd56,6'd57,6'd58,6'd71,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd73: Enemy_img = 4'd14;
//6'd50,6'd53,6'd54,6'd56,6'd57,6'd72,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd58,6'd59,6'd64,6'd65: Enemy_img = 4'd7;
//6'd47,6'd67,6'd68,6'd69,6'd70,6'd76,6'd77: Enemy_img = 4'd14;
//6'd46,6'd56,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd66,6'd67,6'd68,6'd69,6'd76,6'd77: Enemy_img = 4'd14;
//6'd45,6'd46,6'd52,6'd53,6'd54,6'd70,6'd71,6'd73,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd63: Enemy_img = 4'd6;
//6'd49,6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd45,6'd46,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd71,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd51,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd45,6'd46,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd70,6'd72,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd75: Enemy_img = 4'd13;
//6'd47,6'd48,6'd50,6'd51,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd14;
//6'd45,6'd46,6'd52,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd69,6'd71,6'd72,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd60,6'd61,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd56,6'd57,6'd59,6'd60,6'd61,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd57,6'd61,6'd62,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd58,6'd59,6'd61,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd61,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63: Enemy_img = 4'd14;
//6'd60,6'd61,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd14;
//6'd61,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd14;
//6'd61,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd56,6'd59,6'd61,6'd62,6'd64,6'd65,6'd67,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd51,6'd56,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd67: Enemy_img = 4'd14;
//6'd50,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd61,6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd67: Enemy_img = 4'd6;
//6'd47: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd40,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd47,6'd48,6'd68: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd68: Enemy_img = 4'd6;
//6'd45,6'd46,6'd66,6'd67: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd47,6'd48,6'd67: Enemy_img = 4'd6;
//6'd46,6'd49,6'd65,6'd66: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd68: Enemy_img = 4'd6;
//6'd49,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd67,6'd68: Enemy_img = 4'd6;
//6'd44,6'd49,6'd50,6'd64,6'd65,6'd66: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd35,6'd37,6'd38,6'd39,6'd41,6'd42: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd45,6'd46,6'd49,6'd50,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd7;
//6'd52,6'd54,6'd55,6'd57,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//6'd35,6'd37,6'd38,6'd39,6'd42,6'd43,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd45,6'd46,6'd51,6'd64,6'd65,6'd66: Enemy_img = 4'd7;
//6'd53,6'd54,6'd56,6'd58: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd42,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd46,6'd64,6'd65,6'd66: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd50,6'd51,6'd68,6'd69,6'd70: Enemy_img = 4'd6;
//6'd46,6'd48,6'd49,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd41,6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd52,6'd68,6'd69,6'd70: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd65,6'd66,6'd67: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd41,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd52,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd66,6'd67: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd41,6'd44,6'd45,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd52,6'd53,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd67,6'd68,6'd69: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd65: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd62,6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd52,6'd53,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd50,6'd51,6'd68,6'd69,6'd70: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd42,6'd44,6'd45,6'd46,6'd62,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd52,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd50,6'd51,6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd30,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd45,6'd46,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd50,6'd51,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd37,6'd38,6'd42,6'd43,6'd45,6'd46,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd31,6'd32,6'd34,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd75,6'd77,6'd78: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd46,6'd50,6'd51,6'd52,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd7;
//6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd76,6'd77,6'd79,6'd87,6'd89: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd52,6'd66,6'd75,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd6;
//6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd7;
//6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd67,6'd68,6'd71,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd52,6'd63,6'd66,6'd69,6'd70,6'd75,6'd76,6'd82,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33: Enemy_img = 4'd6;
//6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd7;
//6'd48,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd65,6'd69,6'd71,6'd72,6'd73,6'd74,6'd78,6'd83,6'd86: Enemy_img = 4'd14;
//6'd42,6'd49,6'd50,6'd53,6'd64,6'd66,6'd67,6'd68,6'd70,6'd77,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38: Enemy_img = 4'd7;
//6'd48,6'd49,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd79,6'd80,6'd81,6'd85,6'd86: Enemy_img = 4'd14;
//6'd40,6'd43,6'd47,6'd50,6'd53,6'd64,6'd65,6'd70,6'd71,6'd74,6'd75,6'd78,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd87: Enemy_img = 4'd6;
//6'd36,6'd37: Enemy_img = 4'd7;
//6'd47,6'd51,6'd52,6'd55,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd75,6'd76,6'd80,6'd81,6'd84: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd48,6'd49,6'd50,6'd53,6'd54,6'd71,6'd72,6'd73,6'd78,6'd79,6'd82,6'd83,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd6;
//6'd37,6'd38: Enemy_img = 4'd7;
//6'd57: Enemy_img = 4'd9;
//6'd56: Enemy_img = 4'd10;
//6'd48,6'd49,6'd51,6'd52,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd72,6'd75,6'd76,6'd79,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd50,6'd53,6'd69,6'd70,6'd71,6'd73,6'd74,6'd78,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd86,6'd87: Enemy_img = 4'd6;
//6'd37,6'd38: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59: Enemy_img = 4'd9;
//6'd54,6'd55,6'd56: Enemy_img = 4'd10;
//6'd47,6'd48,6'd49,6'd51,6'd61,6'd63,6'd64,6'd65,6'd66,6'd71,6'd72,6'd73,6'd75,6'd76,6'd79,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd45,6'd46,6'd50,6'd67,6'd68,6'd69,6'd70,6'd74,6'd78,6'd80,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd85,6'd86: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55: Enemy_img = 4'd9;
//6'd56: Enemy_img = 4'd10;
//6'd48,6'd49,6'd61,6'd62,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd79,6'd80,6'd82: Enemy_img = 4'd14;
//6'd41,6'd42,6'd47,6'd50,6'd51,6'd66,6'd70,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd86,6'd87: Enemy_img = 4'd6;
//6'd37,6'd38: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd46,6'd50,6'd51,6'd52,6'd53,6'd70,6'd78,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd85,6'd86: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38,6'd84: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd52,6'd71,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd85,6'd86: Enemy_img = 4'd6;
//6'd37,6'd38,6'd83,6'd84: Enemy_img = 4'd7;
//6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd72,6'd74,6'd75,6'd76,6'd79,6'd80: Enemy_img = 4'd14;
//6'd40,6'd42,6'd43,6'd46,6'd47,6'd51,6'd56,6'd71,6'd73,6'd78,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd2;
//6'd34,6'd35,6'd36,6'd85,6'd86: Enemy_img = 4'd6;
//6'd37,6'd38,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd39,6'd40,6'd44,6'd45,6'd47,6'd48,6'd51,6'd72,6'd74,6'd76,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd59,6'd60: Enemy_img = 4'd2;
//6'd34,6'd35,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd36,6'd37,6'd82,6'd83: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd79: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd47,6'd48,6'd50,6'd55,6'd74,6'd75,6'd77,6'd78,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd2;
//6'd33,6'd34,6'd35,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd36,6'd37,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd52,6'd58,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd76: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd44,6'd45,6'd51,6'd53,6'd54,6'd75,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd2;
//6'd33,6'd34,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd35,6'd36,6'd82,6'd83: Enemy_img = 4'd7;
//6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd78: Enemy_img = 4'd14;
//6'd39,6'd42,6'd43,6'd45,6'd46,6'd48,6'd51,6'd52,6'd53,6'd58,6'd74,6'd75,6'd77,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd35,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd53,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd52,6'd54,6'd57,6'd73,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61: Enemy_img = 4'd2;
//6'd32,6'd33,6'd34,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd52,6'd53,6'd56,6'd57,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd51,6'd54,6'd74,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd2;
//6'd32,6'd33,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd34,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd56,6'd57,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd51,6'd55,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd2;
//6'd31,6'd32,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd52,6'd53,6'd56,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd46,6'd47,6'd48,6'd49,6'd51,6'd54,6'd55,6'd59,6'd72,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd2;
//6'd31,6'd32,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd51,6'd52,6'd54,6'd55,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd74: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd53,6'd56,6'd60,6'd70,6'd71,6'd72,6'd73,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd74,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd52,6'd53,6'd55,6'd56,6'd57,6'd60,6'd62,6'd63,6'd64,6'd66,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd36,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd54,6'd58,6'd59,6'd61,6'd67,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd51,6'd53,6'd56,6'd58,6'd60,6'd62,6'd63,6'd65,6'd66,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd31,6'd33,6'd34,6'd36,6'd37,6'd44,6'd46,6'd47,6'd49,6'd50,6'd52,6'd54,6'd55,6'd57,6'd59,6'd61,6'd67,6'd68,6'd72,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd62,6'd63,6'd66,6'd67,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd31,6'd33,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd46,6'd54,6'd56,6'd58,6'd59,6'd60,6'd61,6'd68,6'd72,6'd75,6'd76,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd64,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd66,6'd67,6'd69,6'd70,6'd73,6'd74,6'd78: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd43,6'd44,6'd45,6'd47,6'd57,6'd58,6'd62,6'd68,6'd71,6'd72,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd61,6'd63,6'd64,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd68,6'd69,6'd70,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd59,6'd67,6'd71,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd62,6'd63,6'd64,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd68,6'd69,6'd70,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd27,6'd28,6'd31,6'd33,6'd36,6'd38,6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd55,6'd56,6'd57,6'd67,6'd71,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd65,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd63,6'd64,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd68,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82: Enemy_img = 4'd14;
//6'd41,6'd43,6'd47,6'd48,6'd50,6'd51,6'd52,6'd55,6'd56,6'd58,6'd59,6'd60,6'd67,6'd69,6'd70,6'd71,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd62,6'd63,6'd64,6'd65,6'd66,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd37,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd69,6'd71,6'd72,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd44,6'd47,6'd50,6'd51,6'd54,6'd56,6'd58,6'd59,6'd68,6'd70,6'd73,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd63,6'd64,6'd65,6'd93,6'd94: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd40,6'd66,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd69,6'd71,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd14;
//6'd49,6'd50,6'd53,6'd54,6'd58,6'd59,6'd60,6'd68,6'd70,6'd72,6'd73,6'd75,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd63,6'd64,6'd65,6'd94,6'd96: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd66,6'd67,6'd89,6'd91,6'd92: Enemy_img = 4'd7;
//6'd70,6'd72,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd69,6'd71,6'd73,6'd75,6'd76,6'd82,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd65,6'd66,6'd67: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd64: Enemy_img = 4'd7;
//6'd70,6'd71,6'd76,6'd78,6'd79,6'd80,6'd81,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd93,6'd95: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd60,6'd69,6'd72,6'd73,6'd75,6'd77,6'd82,6'd83,6'd84,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd72,6'd76,6'd79,6'd80,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd53,6'd56,6'd57,6'd58,6'd59,6'd61,6'd69,6'd71,6'd73,6'd75,6'd77,6'd78,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd64,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd67,6'd83: Enemy_img = 4'd7;
//6'd75,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59,6'd61,6'd71,6'd72,6'd73,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd86,6'd87,6'd88,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd65,6'd68,6'd69,6'd78,6'd86: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd66,6'd67,6'd83,6'd84: Enemy_img = 4'd7;
//6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd58,6'd59,6'd60,6'd62,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd81,6'd88,6'd89,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd64,6'd65,6'd78,6'd79,6'd81,6'd86: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd66,6'd67,6'd68,6'd69,6'd70,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd89,6'd90,6'd91,6'd93: Enemy_img = 4'd14;
//6'd52,6'd60,6'd61,6'd72,6'd73,6'd75,6'd76,6'd88,6'd92,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd65,6'd78,6'd80,6'd81,6'd82,6'd83,6'd85: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd66,6'd67,6'd68,6'd69,6'd70,6'd79,6'd84: Enemy_img = 4'd7;
//6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd61,6'd72,6'd74,6'd75,6'd76,6'd87,6'd88,6'd89,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd77,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd51,6'd53,6'd54,6'd55,6'd56,6'd62,6'd73,6'd75,6'd87,6'd88,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd76,6'd77,6'd85: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd88,6'd89,6'd91: Enemy_img = 4'd14;
//6'd54,6'd57,6'd58,6'd86,6'd87,6'd90,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd52,6'd55,6'd57,6'd58,6'd83,6'd84,6'd86,6'd87,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd73,6'd75: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd84,6'd87,6'd88: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd55,6'd56,6'd60,6'd83,6'd85,6'd86,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd72,6'd73: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd81: Enemy_img = 4'd7;
//6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd56,6'd77,6'd78,6'd79,6'd82,6'd83,6'd86,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd58,6'd59,6'd66,6'd72,6'd73: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd7;
//6'd83,6'd84: Enemy_img = 4'd14;
//6'd51,6'd52,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd70,6'd71,6'd73: Enemy_img = 4'd7;
//6'd77,6'd80,6'd83,6'd85,6'd86: Enemy_img = 4'd14;
//6'd51,6'd52,6'd74,6'd75,6'd76,6'd78,6'd79,6'd81,6'd82,6'd84,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd59,6'd66,6'd67,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd78,6'd80,6'd81,6'd82,6'd83,6'd85: Enemy_img = 4'd14;
//6'd51,6'd52,6'd74,6'd76,6'd77,6'd79,6'd84,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd58,6'd63,6'd71: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd54,6'd59,6'd60,6'd61,6'd62,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd7;
//6'd75,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd14;
//6'd50,6'd74,6'd78,6'd79,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd57,6'd58,6'd71,6'd72: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd74,6'd75,6'd76,6'd78,6'd83,6'd84,6'd88: Enemy_img = 4'd14;
//6'd81,6'd82,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd57,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd84,6'd88,6'd89: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd82,6'd83,6'd85,6'd86,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd53,6'd54,6'd55,6'd57,6'd73: Enemy_img = 4'd6;
//6'd46,6'd56,6'd59,6'd60,6'd61,6'd72: Enemy_img = 4'd7;
//6'd87: Enemy_img = 4'd13;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd88,6'd89: Enemy_img = 4'd14;
//6'd49,6'd50,6'd65,6'd66,6'd69,6'd70,6'd84,6'd85,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd54,6'd55,6'd56,6'd72: Enemy_img = 4'd6;
//6'd45,6'd46,6'd61,6'd73: Enemy_img = 4'd7;
//6'd87: Enemy_img = 4'd13;
//6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd65,6'd66,6'd70,6'd83,6'd85,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd56,6'd73,6'd74: Enemy_img = 4'd6;
//6'd75,6'd76: Enemy_img = 4'd7;
//6'd88: Enemy_img = 4'd13;
//6'd79,6'd80,6'd81,6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd14;
//6'd47,6'd49,6'd64,6'd65,6'd68,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd73,6'd74: Enemy_img = 4'd6;
//6'd72,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd88: Enemy_img = 4'd13;
//6'd79,6'd80,6'd81,6'd82,6'd83,6'd86,6'd87: Enemy_img = 4'd14;
//6'd46,6'd47,6'd51,6'd52,6'd53,6'd60,6'd63,6'd64,6'd68,6'd69,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd71,6'd72: Enemy_img = 4'd7;
//6'd79,6'd80,6'd81,6'd82,6'd86: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd55,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd76: Enemy_img = 4'd6;
//6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd7;
//6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd68,6'd69,6'd70,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73,6'd76: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd43,6'd45,6'd47,6'd49,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd63,6'd64,6'd66,6'd67,6'd69,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd43,6'd44,6'd62,6'd63,6'd71,6'd72,6'd75,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd42,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd60,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd77,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd13;
//6'd61,6'd62,6'd64,6'd65,6'd66,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd59,6'd60,6'd67,6'd72,6'd74,6'd76,6'd77,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd65,6'd66,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd71,6'd72,6'd75,6'd77,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd13;
//6'd62,6'd63,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd60,6'd61,6'd74,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd14;
//6'd60,6'd61,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd14;
//6'd77,6'd78,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd14;
//6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd14;
//6'd50,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd46,6'd48,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd45,6'd46,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd43,6'd45,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd40,6'd42,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54: Enemy_img = 4'd6;
//6'd52: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54: Enemy_img = 4'd6;
//6'd52: Enemy_img = 4'd7;
//6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd37,6'd39,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53: Enemy_img = 4'd7;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd33,6'd35: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd33,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd70,6'd73: Enemy_img = 4'd6;
//6'd32,6'd33,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd79: Enemy_img = 4'd14;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd35,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd51,6'd77,6'd78: Enemy_img = 4'd14;
//6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd35,6'd36,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd6;
//6'd33,6'd34,6'd37,6'd38,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd7;
//6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//6'd27,6'd28,6'd51,6'd52,6'd76,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd70,6'd74,6'd75,6'd77: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd52,6'd53,6'd72,6'd73,6'd76,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd79: Enemy_img = 4'd6;
//6'd33,6'd39,6'd40,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd57,6'd68,6'd69,6'd70,6'd71,6'd76,6'd77: Enemy_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd52,6'd53,6'd72,6'd73,6'd74,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd67,6'd69,6'd70,6'd73,6'd76: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd53,6'd59,6'd66,6'd68,6'd71,6'd72,6'd74,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd79: Enemy_img = 4'd6;
//6'd34,6'd35,6'd39: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd72,6'd73,6'd76: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd52,6'd59,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd42,6'd43,6'd79,6'd80: Enemy_img = 4'd6;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd72,6'd75: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd58,6'd71,6'd73,6'd74,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd43,6'd44,6'd79,6'd80: Enemy_img = 4'd6;
//6'd36,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32,6'd33,6'd34,6'd57,6'd58,6'd61,6'd62,6'd67,6'd71,6'd73,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd43,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd7;
//6'd46,6'd50,6'd52,6'd53,6'd56,6'd57,6'd61,6'd62,6'd64,6'd65,6'd67,6'd68,6'd69,6'd73,6'd75: Enemy_img = 4'd14;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd58,6'd59,6'd60,6'd63,6'd66,6'd71,6'd72,6'd74,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd43,6'd44,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd78: Enemy_img = 4'd7;
//6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd66,6'd68,6'd69,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd56,6'd59,6'd64,6'd65,6'd67,6'd70,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd78: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd73,6'd74: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd32,6'd33,6'd35,6'd36,6'd37,6'd56,6'd57,6'd58,6'd64,6'd68,6'd69,6'd70,6'd72,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd42,6'd80,6'd81: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd73,6'd74: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd30,6'd31,6'd34,6'd36,6'd37,6'd38,6'd57,6'd63,6'd69,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd77,6'd78: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd37,6'd38,6'd39,6'd40,6'd43,6'd44,6'd62,6'd64,6'd72,6'd73,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd78,6'd79: Enemy_img = 4'd7;
//6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36,6'd38,6'd39,6'd40,6'd42,6'd43,6'd45,6'd61,6'd65,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd55,6'd57,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd70,6'd74: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd39,6'd46,6'd60,6'd66,6'd68,6'd69,6'd71,6'd73,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd52,6'd53: Enemy_img = 4'd9;
//6'd44,6'd45,6'd46,6'd48,6'd49,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd71,6'd72,6'd74: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd42,6'd43,6'd47,6'd67,6'd68,6'd70,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd52,6'd54: Enemy_img = 4'd9;
//6'd51: Enemy_img = 4'd10;
//6'd42,6'd43,6'd45,6'd46,6'd47,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd30,6'd31,6'd33,6'd35,6'd36,6'd37,6'd38,6'd44,6'd48,6'd71,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd50,6'd51: Enemy_img = 4'd10;
//6'd43,6'd45,6'd46,6'd47,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd66,6'd67,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd25,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd44,6'd71,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd49,6'd50: Enemy_img = 4'd9;
//6'd42,6'd46,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd20,6'd21,6'd33,6'd34,6'd35,6'd36,6'd43,6'd44,6'd45,6'd70,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd48: Enemy_img = 4'd9;
//6'd43,6'd44,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd34,6'd38,6'd41,6'd42,6'd45,6'd46,6'd49,6'd71,6'd73,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd24,6'd25,6'd26,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd53,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd46,6'd47,6'd48,6'd52,6'd71,6'd72,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd2;
//6'd25,6'd26,6'd27,6'd28,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd40,6'd42,6'd43,6'd45,6'd46,6'd49,6'd70,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd47,6'd71,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54: Enemy_img = 4'd2;
//6'd28,6'd29,6'd30,6'd31,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd49,6'd50,6'd51,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd52,6'd53,6'd55,6'd56,6'd69,6'd71,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd58,6'd61: Enemy_img = 4'd2;
//6'd29,6'd30,6'd31,6'd32,6'd91,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92: Enemy_img = 4'd7;
//6'd49,6'd50,6'd63,6'd64,6'd65,6'd67,6'd71,6'd72,6'd73,6'd74,6'd99,6'd101: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd51,6'd52,6'd55,6'd56,6'd75,6'd76,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd2;
//6'd30,6'd31,6'd32: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd56,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd73,6'd74,6'd78,6'd79,6'd80,6'd97,6'd100: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd71,6'd72,6'd75,6'd76,6'd77,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33: Enemy_img = 4'd6;
//6'd34,6'd35,6'd85,6'd86,6'd88,6'd89,6'd91: Enemy_img = 4'd7;
//6'd51,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd68,6'd69,6'd70,6'd71,6'd74,6'd78,6'd79,6'd80,6'd81,6'd83,6'd94,6'd95,6'd96,6'd97,6'd99: Enemy_img = 4'd14;
//6'd37,6'd40,6'd42,6'd43,6'd45,6'd50,6'd52,6'd53,6'd59,6'd67,6'd72,6'd73,6'd75,6'd77,6'd98,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd31,6'd32,6'd33: Enemy_img = 4'd6;
//6'd34,6'd35: Enemy_img = 4'd7;
//6'd51,6'd52,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd38,6'd42,6'd43,6'd44,6'd47,6'd53,6'd54,6'd59,6'd60,6'd68,6'd72,6'd73,6'd75,6'd77,6'd85,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd2;
//6'd32,6'd33,6'd34: Enemy_img = 4'd6;
//6'd35,6'd36: Enemy_img = 4'd7;
//6'd52,6'd53,6'd56,6'd59,6'd62,6'd63,6'd66,6'd67,6'd68,6'd70,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd54,6'd55,6'd60,6'd61,6'd69,6'd71,6'd72,6'd75,6'd76,6'd77,6'd86,6'd90,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd6;
//6'd35,6'd36: Enemy_img = 4'd7;
//6'd52,6'd55,6'd60,6'd63,6'd67,6'd68,6'd70,6'd71,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd88,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd38,6'd39,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd51,6'd53,6'd54,6'd56,6'd59,6'd61,6'd62,6'd69,6'd72,6'd73,6'd75,6'd76,6'd77,6'd84,6'd86,6'd87,6'd89,6'd90,6'd91,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34: Enemy_img = 4'd6;
//6'd35,6'd36,6'd65: Enemy_img = 4'd7;
//6'd52,6'd53,6'd56,6'd57,6'd58,6'd61,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd38,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd51,6'd54,6'd55,6'd59,6'd60,6'd62,6'd68,6'd73,6'd74,6'd75,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd89: Enemy_img = 4'd6;
//6'd35,6'd36,6'd65,6'd66,6'd88: Enemy_img = 4'd7;
//6'd52,6'd54,6'd56,6'd57,6'd59,6'd70,6'd74,6'd80,6'd81,6'd82,6'd83,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd51,6'd53,6'd55,6'd58,6'd60,6'd63,6'd69,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd84,6'd85,6'd91,6'd92,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd67,6'd90: Enemy_img = 4'd6;
//6'd35,6'd63,6'd64,6'd65,6'd66,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd71,6'd72,6'd78,6'd79,6'd82,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd56,6'd57,6'd58,6'd70,6'd73,6'd74,6'd75,6'd76,6'd80,6'd81,6'd83,6'd84,6'd85,6'd91,6'd92,6'd93,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd68,6'd89,6'd90: Enemy_img = 4'd6;
//6'd35,6'd64,6'd65,6'd66,6'd67,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd52,6'd72,6'd73,6'd75,6'd79,6'd93,6'd94: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd71,6'd74,6'd76,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd92,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd65,6'd67,6'd68,6'd82,6'd85,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd66,6'd69,6'd87: Enemy_img = 4'd7;
//6'd73,6'd74,6'd75,6'd79,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd37,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd53,6'd59,6'd60,6'd62,6'd72,6'd76,6'd80,6'd81,6'd92,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd66,6'd67,6'd68,6'd69,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd35,6'd70: Enemy_img = 4'd7;
//6'd76,6'd93,6'd94: Enemy_img = 4'd14;
//6'd36,6'd40,6'd41,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd56,6'd58,6'd59,6'd61,6'd62,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd91,6'd92,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd68,6'd69,6'd70,6'd71,6'd73,6'd82,6'd83: Enemy_img = 4'd6;
//6'd67,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd93,6'd94: Enemy_img = 4'd14;
//6'd36,6'd37,6'd40,6'd43,6'd44,6'd46,6'd48,6'd52,6'd53,6'd54,6'd55,6'd58,6'd59,6'd61,6'd62,6'd63,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd90,6'd91,6'd92,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd82: Enemy_img = 4'd6;
//6'd68,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd93,6'd94: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd45,6'd46,6'd47,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd62,6'd63,6'd64,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd89,6'd90,6'd91,6'd92,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd69,6'd70,6'd73,6'd74,6'd82,6'd83: Enemy_img = 4'd6;
//6'd71,6'd72,6'd75,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd90,6'd91: Enemy_img = 4'd14;
//6'd36,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd57,6'd58,6'd61,6'd62,6'd64,6'd65,6'd77,6'd78,6'd80,6'd88,6'd89,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd70,6'd82,6'd83: Enemy_img = 4'd6;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd81,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd90,6'd93: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd40,6'd42,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd57,6'd58,6'd59,6'd61,6'd63,6'd65,6'd66,6'd78,6'd79,6'd88,6'd89,6'd91,6'd92,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd69,6'd70,6'd71,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd92: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd44,6'd46,6'd51,6'd54,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd87,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd79,6'd80: Enemy_img = 4'd6;
//6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81: Enemy_img = 4'd7;
//6'd90,6'd93,6'd96: Enemy_img = 4'd14;
//6'd34,6'd36,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd53,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd91,6'd92,6'd94,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80: Enemy_img = 4'd6;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd87,6'd88,6'd89,6'd90,6'd93,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd66,6'd67,6'd83,6'd84,6'd85,6'd86,6'd91,6'd92,6'd94,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd6;
//6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81: Enemy_img = 4'd7;
//6'd84,6'd85,6'd88,6'd89,6'd92,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd34,6'd37,6'd38,6'd40,6'd68,6'd82,6'd83,6'd86,6'd87,6'd90,6'd91,6'd93,6'd94,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd6;
//6'd44,6'd45,6'd47,6'd48,6'd50,6'd51,6'd52,6'd54,6'd55,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81: Enemy_img = 4'd7;
//6'd96: Enemy_img = 4'd13;
//6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd80: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd97: Enemy_img = 4'd13;
//6'd85,6'd95,6'd96,6'd98: Enemy_img = 4'd14;
//6'd33,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd82,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd74,6'd76,6'd77,6'd80: Enemy_img = 4'd6;
//6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd75,6'd78,6'd79: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd96,6'd97: Enemy_img = 4'd14;
//6'd32,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd82,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd81: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd96: Enemy_img = 4'd14;
//6'd58,6'd61,6'd63,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd73,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd72,6'd74,6'd76,6'd77: Enemy_img = 4'd7;
//6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd63,6'd64,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd83: Enemy_img = 4'd6;
//6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd81,6'd82: Enemy_img = 4'd7;
//6'd85,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd68,6'd69,6'd71,6'd72,6'd82,6'd83: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd70,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62,6'd79,6'd80,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd68,6'd83,6'd84,6'd85,6'd86,6'd88: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd69,6'd70,6'd71,6'd72,6'd87: Enemy_img = 4'd7;
//6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd60,6'd61,6'd76,6'd80,6'd81,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd67,6'd68,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd69,6'd70,6'd71,6'd72,6'd83: Enemy_img = 4'd7;
//6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd75,6'd76,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd67,6'd68,6'd84,6'd85,6'd88: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd66,6'd69,6'd70,6'd71,6'd72,6'd83,6'd86: Enemy_img = 4'd7;
//6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd60,6'd61,6'd75,6'd76,6'd79,6'd80,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd68,6'd85: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd83,6'd84: Enemy_img = 4'd7;
//6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd61,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd67,6'd68,6'd84,6'd86: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd64,6'd65,6'd66,6'd83: Enemy_img = 4'd7;
//6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd60,6'd75,6'd76,6'd79,6'd80,6'd81,6'd87,6'd88,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd64,6'd66,6'd67,6'd68: Enemy_img = 4'd6;
//6'd57,6'd58,6'd59,6'd65: Enemy_img = 4'd7;
//6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd62,6'd75,6'd76,6'd81,6'd84,6'd87,6'd88,6'd89,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd6;
//6'd57,6'd58: Enemy_img = 4'd7;
//6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd61,6'd72,6'd73,6'd75,6'd79,6'd83,6'd84,6'd85,6'd88,6'd89,6'd90,6'd91,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd6;
//6'd58,6'd59: Enemy_img = 4'd7;
//6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//6'd60,6'd61,6'd71,6'd73,6'd74,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88,6'd90,6'd91,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd6;
//6'd57,6'd58: Enemy_img = 4'd7;
//6'd93,6'd94: Enemy_img = 4'd14;
//6'd60,6'd61,6'd62,6'd71,6'd72,6'd74,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83,6'd84,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd6;
//6'd58: Enemy_img = 4'd7;
//6'd94: Enemy_img = 4'd14;
//6'd61,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd79,6'd81,6'd82,6'd86,6'd87,6'd89,6'd91,6'd92,6'd93,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57: Enemy_img = 4'd6;
//6'd95: Enemy_img = 4'd14;
//6'd59,6'd60,6'd62,6'd65,6'd68,6'd69,6'd70,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57: Enemy_img = 4'd6;
//6'd78: Enemy_img = 4'd13;
//6'd75,6'd80: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd67,6'd81,6'd94,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd79: Enemy_img = 4'd13;
//6'd75,6'd76,6'd77,6'd80: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57: Enemy_img = 4'd6;
//6'd79: Enemy_img = 4'd13;
//6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd58,6'd61,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78: Enemy_img = 4'd14;
//6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd59,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43: Enemy_img = 4'd14;
//6'd41,6'd42,6'd44: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd39,6'd40: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd38,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd6;
//6'd45: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd37,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd6;
//6'd45: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd35,6'd36,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd45,6'd46: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd72: Enemy_img = 4'd14;
//6'd34,6'd35,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd67,6'd68: Enemy_img = 4'd6;
//6'd45,6'd46: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd33,6'd43: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd71: Enemy_img = 4'd14;
//6'd32,6'd43,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd7;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd68,6'd69,6'd71: Enemy_img = 4'd14;
//6'd30,6'd31,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd74: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd68,6'd69,6'd71: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd66,6'd67,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd74: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd65,6'd66,6'd71: Enemy_img = 4'd14;
//6'd27,6'd28,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd63,6'd64,6'd65,6'd67,6'd68,6'd71: Enemy_img = 4'd14;
//6'd66,6'd69,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd43,6'd44,6'd45,6'd46,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71: Enemy_img = 4'd14;
//6'd61,6'd66,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd67,6'd68,6'd70,6'd71: Enemy_img = 4'd14;
//6'd47,6'd48,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd28,6'd31: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd67,6'd68: Enemy_img = 4'd14;
//6'd48,6'd66,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd27,6'd28,6'd29,6'd32,6'd74: Enemy_img = 4'd7;
//6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd68,6'd69: Enemy_img = 4'd14;
//6'd48,6'd54,6'd63,6'd67,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd27,6'd28,6'd29,6'd32,6'd33,6'd34,6'd74: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd48,6'd54,6'd57,6'd58,6'd62,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd74,6'd75: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd64,6'd65,6'd69,6'd70: Enemy_img = 4'd14;
//6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd74,6'd75: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd52,6'd53,6'd54,6'd57,6'd58,6'd59,6'd62,6'd63,6'd66,6'd67,6'd70,6'd71: Enemy_img = 4'd14;
//6'd23,6'd24,6'd55,6'd56,6'd60,6'd61,6'd64,6'd65,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd55,6'd56,6'd60,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd39,6'd40,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd38,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd52,6'd56,6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd70,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd39,6'd40,6'd41,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd31,6'd32,6'd35,6'd36,6'd37,6'd38,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd71: Enemy_img = 4'd14;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd54,6'd59,6'd61,6'd62,6'd68,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd40,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd33,6'd36,6'd37,6'd38,6'd39,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd69: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd58,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd40,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd38,6'd39,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd70: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd58,6'd64,6'd68,6'd69,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd99: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd32,6'd33,6'd34,6'd68,6'd69,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd67,6'd70,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd21,6'd22,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd41,6'd42,6'd43,6'd68,6'd69,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90,6'd93: Enemy_img = 4'd6;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd91,6'd92: Enemy_img = 4'd7;
//6'd50,6'd51: Enemy_img = 4'd9;
//6'd42,6'd45,6'd46,6'd47,6'd48,6'd54,6'd55,6'd56,6'd57,6'd64,6'd65,6'd67,6'd68,6'd96,6'd98: Enemy_img = 4'd14;
//6'd22,6'd23,6'd24,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd43,6'd44,6'd69,6'd70,6'd71,6'd74,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52: Enemy_img = 4'd9;
//6'd49: Enemy_img = 4'd10;
//6'd42,6'd43,6'd44,6'd47,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd71,6'd72,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd32,6'd36,6'd37,6'd38,6'd41,6'd45,6'd46,6'd69,6'd70,6'd74,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd50: Enemy_img = 4'd9;
//6'd49: Enemy_img = 4'd10;
//6'd43,6'd44,6'd45,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd37,6'd38,6'd41,6'd42,6'd46,6'd69,6'd72,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd48,6'd49: Enemy_img = 4'd10;
//6'd41,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd40,6'd42,6'd43,6'd46,6'd70,6'd71,6'd74,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49: Enemy_img = 4'd9;
//6'd41,6'd42,6'd44,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd72,6'd73,6'd78,6'd79,6'd80,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd43,6'd69,6'd74,6'd75,6'd77,6'd89,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56: Enemy_img = 4'd2;
//6'd41,6'd50,6'd51,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67,6'd70,6'd71,6'd72,6'd73,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd40,6'd42,6'd43,6'd44,6'd45,6'd48,6'd52,6'd68,6'd74,6'd75,6'd77,6'd84,6'd85,6'd89,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd2;
//6'd43,6'd44,6'd50,6'd51,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd69,6'd70,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd42,6'd45,6'd46,6'd48,6'd71,6'd72,6'd75,6'd77,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd60: Enemy_img = 4'd2;
//6'd41,6'd42,6'd43,6'd44,6'd50,6'd51,6'd56,6'd57,6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd33,6'd34,6'd37,6'd38,6'd40,6'd45,6'd46,6'd55,6'd72,6'd75,6'd77,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd92,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd58,6'd59: Enemy_img = 4'd2;
//6'd89,6'd90: Enemy_img = 4'd6;
//6'd28,6'd29,6'd30,6'd31,6'd87: Enemy_img = 4'd7;
//6'd41,6'd49,6'd50,6'd51,6'd62,6'd63,6'd64,6'd66,6'd69,6'd70,6'd71,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd94: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd36,6'd37,6'd38,6'd40,6'd42,6'd47,6'd52,6'd55,6'd56,6'd67,6'd68,6'd72,6'd75,6'd76,6'd84,6'd85,6'd92,6'd93,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd57,6'd58: Enemy_img = 4'd2;
//6'd90: Enemy_img = 4'd6;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd49,6'd50,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd70,6'd71,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd94,6'd95: Enemy_img = 4'd14;
//6'd20,6'd21,6'd22,6'd35,6'd36,6'd37,6'd38,6'd48,6'd51,6'd52,6'd68,6'd69,6'd72,6'd73,6'd76,6'd85,6'd92,6'd93,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd2;
//6'd90: Enemy_img = 4'd6;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd82,6'd94,6'd95: Enemy_img = 4'd14;
//6'd20,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd59,6'd60,6'd69,6'd74,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd92,6'd93,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd2;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd7;
//6'd51,6'd52,6'd55,6'd56,6'd60,6'd62,6'd63,6'd64,6'd68,6'd70,6'd71,6'd72,6'd75,6'd79,6'd80,6'd94,6'd95: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd53,6'd54,6'd61,6'd69,6'd73,6'd74,6'd76,6'd81,6'd82,6'd83,6'd84,6'd93,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd66,6'd67: Enemy_img = 4'd7;
//6'd52,6'd53,6'd56,6'd60,6'd61,6'd64,6'd76,6'd80,6'd94,6'd95: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd46,6'd51,6'd54,6'd55,6'd62,6'd63,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd79,6'd81,6'd93,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd68,6'd83,6'd84: Enemy_img = 4'd6;
//6'd34,6'd35,6'd36,6'd66,6'd67,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd62,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd40,6'd41,6'd43,6'd44,6'd48,6'd51,6'd55,6'd57,6'd60,6'd61,6'd63,6'd64,6'd71,6'd72,6'd77,6'd78,6'd80,6'd81,6'd82,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd69,6'd70,6'd84: Enemy_img = 4'd6;
//6'd34,6'd35,6'd36,6'd64,6'd65,6'd66,6'd67,6'd68,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd53,6'd54,6'd58,6'd59,6'd60,6'd75,6'd76,6'd77,6'd92,6'd93: Enemy_img = 4'd14;
//6'd38,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd55,6'd56,6'd57,6'd61,6'd73,6'd74,6'd78,6'd80,6'd81,6'd82,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd32,6'd33,6'd34,6'd68,6'd69,6'd70,6'd84: Enemy_img = 4'd6;
//6'd35,6'd36,6'd37,6'd65,6'd66,6'd67,6'd71,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd53,6'd58,6'd92,6'd94,6'd95: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd57,6'd59,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd90,6'd91,6'd93,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd84,6'd85: Enemy_img = 4'd6;
//6'd36,6'd37,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd55,6'd56,6'd92,6'd95,6'd98,6'd99: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd57,6'd58,6'd61,6'd62,6'd78,6'd79,6'd80,6'd82,6'd91,6'd93,6'd94,6'd96,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd33,6'd34,6'd35,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd85: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38,6'd84: Enemy_img = 4'd7;
//6'd54,6'd55,6'd92,6'd93,6'd95,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd53,6'd56,6'd57,6'd61,6'd62,6'd64,6'd79,6'd80,6'd89,6'd90,6'd91,6'd94,6'd96,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd71,6'd72,6'd73,6'd83,6'd84: Enemy_img = 4'd6;
//6'd37,6'd38,6'd70,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd92,6'd93,6'd95,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd61,6'd64,6'd65,6'd81,6'd87,6'd88,6'd89,6'd90,6'd91,6'd94,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd71,6'd72,6'd73,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd37,6'd38,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd99,6'd100: Enemy_img = 4'd13;
//6'd90,6'd91,6'd92,6'd94,6'd95,6'd96,6'd101: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd58,6'd61,6'd64,6'd65,6'd66,6'd67,6'd86,6'd87,6'd88,6'd89,6'd93,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd72,6'd73,6'd82,6'd83: Enemy_img = 4'd6;
//6'd37,6'd38,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84: Enemy_img = 4'd7;
//6'd101: Enemy_img = 4'd13;
//6'd88,6'd89,6'd99,6'd100: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd56,6'd57,6'd58,6'd62,6'd64,6'd67,6'd68,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd73,6'd74,6'd83: Enemy_img = 4'd6;
//6'd37,6'd38,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84: Enemy_img = 4'd7;
//6'd88,6'd99,6'd100: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd64,6'd66,6'd85,6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd74,6'd83: Enemy_img = 4'd6;
//6'd38,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84: Enemy_img = 4'd7;
//6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd40,6'd42,6'd43,6'd46,6'd47,6'd49,6'd53,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd86,6'd96,6'd97,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd83,6'd84: Enemy_img = 4'd6;
//6'd38,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd39,6'd40,6'd43,6'd44,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd86,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd84: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd60,6'd61,6'd62,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd80,6'd81,6'd82,6'd84: Enemy_img = 4'd6;
//6'd78,6'd79,6'd83,6'd85: Enemy_img = 4'd7;
//6'd88,6'd89,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd39,6'd40,6'd57,6'd60,6'd61: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd92: Enemy_img = 4'd7;
//6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd78,6'd87: Enemy_img = 4'd6;
//6'd79,6'd80,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd39,6'd40,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd78,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd77: Enemy_img = 4'd7;
//6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd84,6'd85,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd74,6'd75,6'd76,6'd77,6'd78,6'd89,6'd90,6'd91,6'd93: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd88,6'd92: Enemy_img = 4'd7;
//6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd63,6'd64,6'd65,6'd66,6'd68,6'd84,6'd85,6'd86,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd72,6'd73,6'd74,6'd75,6'd77,6'd90: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd76,6'd88,6'd89,6'd91: Enemy_img = 4'd7;
//6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd39,6'd42,6'd43,6'd44,6'd63,6'd68,6'd69,6'd81,6'd82,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd90,6'd91: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd74,6'd75,6'd76,6'd77,6'd88,6'd89: Enemy_img = 4'd7;
//6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd39,6'd40,6'd42,6'd65,6'd66,6'd67,6'd70,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd93,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd49,6'd50,6'd51,6'd53,6'd54,6'd73: Enemy_img = 4'd6;
//6'd47,6'd48,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd74,6'd75,6'd76,6'd77,6'd78,6'd89: Enemy_img = 4'd7;
//6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd65,6'd66,6'd67,6'd70,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd93,6'd94,6'd95,6'd96,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd73: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd98,6'd99,6'd100: Enemy_img = 4'd14;
//6'd38,6'd39,6'd66,6'd67,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd73,6'd74: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd71,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd99,6'd100: Enemy_img = 4'd14;
//6'd38,6'd66,6'd67,6'd81,6'd82,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95,6'd97,6'd98,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd74: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd100,6'd101: Enemy_img = 4'd14;
//6'd38,6'd66,6'd67,6'd68,6'd81,6'd82,6'd85,6'd86,6'd89,6'd90,6'd91,6'd96,6'd98,6'd99,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd74: Enemy_img = 4'd6;
//6'd62,6'd63,6'd64,6'd65,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd67,6'd79,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd7;
//6'd67,6'd79,6'd80,6'd83,6'd86,6'd87,6'd88,6'd89,6'd90,6'd93,6'd94,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd62,6'd72,6'd73: Enemy_img = 4'd6;
//6'd63,6'd64,6'd65: Enemy_img = 4'd7;
//6'd68,6'd78,6'd81,6'd82,6'd83,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66: Enemy_img = 4'd7;
//6'd68,6'd78,6'd79,6'd81,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66: Enemy_img = 4'd7;
//6'd87,6'd88: Enemy_img = 4'd14;
//6'd68,6'd69,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64: Enemy_img = 4'd6;
//6'd65,6'd66: Enemy_img = 4'd7;
//6'd86: Enemy_img = 4'd13;
//6'd83,6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd68,6'd69,6'd71,6'd72,6'd73,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64: Enemy_img = 4'd6;
//6'd65,6'd66: Enemy_img = 4'd7;
//6'd87: Enemy_img = 4'd13;
//6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd72,6'd73,6'd75,6'd76,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64: Enemy_img = 4'd6;
//6'd65: Enemy_img = 4'd7;
//6'd85,6'd86: Enemy_img = 4'd14;
//6'd70,6'd73,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65: Enemy_img = 4'd6;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65: Enemy_img = 4'd6;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65: Enemy_img = 4'd6;
//6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd14;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd14;
//6'd63,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd63,6'd81: Enemy_img = 4'd14;
//6'd62,6'd64,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd62,6'd63,6'd65,6'd66,6'd67,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61: Enemy_img = 4'd6;
//6'd82: Enemy_img = 4'd13;
//6'd62,6'd63,6'd64,6'd65,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd14;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81: Enemy_img = 4'd13;
//6'd63,6'd64,6'd65,6'd66,6'd69,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd67,6'd68,6'd70,6'd71,6'd72,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61: Enemy_img = 4'd6;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd79,6'd82,6'd98: Enemy_img = 4'd14;
//6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd84,6'd85,6'd94,6'd95,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61: Enemy_img = 4'd6;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd91,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd89,6'd90,6'd92,6'd93,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61: Enemy_img = 4'd6;
//6'd62: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd78,6'd79,6'd85,6'd86,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd69,6'd75,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd77,6'd80,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd81,6'd84,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61: Enemy_img = 4'd6;
//6'd62,6'd63: Enemy_img = 4'd7;
//6'd64,6'd65,6'd75,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd75,6'd76,6'd78,6'd79,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd65,6'd66,6'd67,6'd73,6'd74,6'd77,6'd80,6'd81,6'd94,6'd95,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd60,6'd68,6'd70,6'd71,6'd72: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63,6'd69: Enemy_img = 4'd7;
//6'd64,6'd65,6'd79,6'd80,6'd83,6'd84,6'd85,6'd87,6'd88,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd66,6'd67,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd93,6'd94,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd71,6'd72,6'd88,6'd90: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd63,6'd68,6'd69,6'd70,6'd87: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd79,6'd80,6'd83,6'd84,6'd85,6'd91: Enemy_img = 4'd14;
//6'd67,6'd75,6'd76,6'd78,6'd81,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd72,6'd89: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd87,6'd88: Enemy_img = 4'd7;
//6'd65,6'd79,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd66,6'd67,6'd77,6'd78,6'd80,6'd81,6'd92,6'd93,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd58,6'd71,6'd72,6'd88,6'd89,6'd92: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd70,6'd73,6'd74,6'd75,6'd76,6'd87,6'd90: Enemy_img = 4'd7;
//6'd64,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd65,6'd66,6'd67,6'd78,6'd79,6'd80,6'd81,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd71,6'd72,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd63,6'd73,6'd74,6'd75,6'd76,6'd87: Enemy_img = 4'd7;
//6'd65,6'd66,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd64,6'd67,6'd68,6'd69,6'd70,6'd78,6'd79,6'd81,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd72,6'd88,6'd89,6'd90,6'd92: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd87,6'd91: Enemy_img = 4'd7;
//6'd64,6'd65,6'd67,6'd80,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd66,6'd68,6'd69,6'd70,6'd78,6'd79,6'd81,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd72,6'd73,6'd75,6'd76,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd74,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd83,6'd84: Enemy_img = 4'd14;
//6'd69,6'd70,6'd79,6'd80,6'd81,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd85,6'd87: Enemy_img = 4'd6;
//6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd86: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd14;
//6'd70,6'd80,6'd81,6'd82,6'd83,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd77,6'd85: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd76,6'd78,6'd80,6'd81,6'd84,6'd86: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd69,6'd70,6'd71,6'd73,6'd74,6'd88,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd7;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd99,6'd100: Enemy_img = 4'd14;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd87,6'd88,6'd90,6'd91,6'd92,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd78,6'd80,6'd81,6'd84: Enemy_img = 4'd6;
//6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd79,6'd82,6'd83: Enemy_img = 4'd7;
//6'd100,6'd101: Enemy_img = 4'd13;
//6'd36,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71: Enemy_img = 4'd14;
//6'd38,6'd68,6'd72,6'd73,6'd74,6'd76,6'd87,6'd90,6'd91,6'd92,6'd94,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd84: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd99,6'd100: Enemy_img = 4'd13;
//6'd37,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd101,6'd102: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd61,6'd68,6'd70,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd100,6'd101,6'd102: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd72,6'd73,6'd74,6'd75,6'd91,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd6;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd44,6'd72,6'd100,6'd101: Enemy_img = 4'd14;
//6'd38,6'd39,6'd43,6'd45,6'd46,6'd48,6'd49,6'd51,6'd52,6'd55,6'd56,6'd58,6'd61,6'd62,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd96,6'd102,6'd103,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd38,6'd39,6'd43,6'd44,6'd45,6'd70,6'd71,6'd99,6'd100: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd83,6'd84: Enemy_img = 4'd6;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd85: Enemy_img = 4'd7;
//6'd38,6'd39,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd71: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd45,6'd53,6'd55,6'd67,6'd69,6'd70,6'd72,6'd95,6'd96,6'd97,6'd100,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd73,6'd74,6'd75,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd41,6'd42,6'd45,6'd46,6'd47,6'd48,6'd50,6'd55,6'd57,6'd58,6'd61,6'd62,6'd65,6'd70,6'd71: Enemy_img = 4'd14;
//6'd39,6'd40,6'd43,6'd44,6'd49,6'd51,6'd56,6'd59,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd72,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd74,6'd86,6'd87: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd85,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd61,6'd67,6'd69,6'd70: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd45,6'd47,6'd49,6'd57,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd71,6'd94,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd73,6'd74,6'd77,6'd78,6'd86,6'd87: Enemy_img = 4'd6;
//6'd75,6'd76,6'd79,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd40,6'd49,6'd50,6'd52,6'd55,6'd58,6'd61,6'd63,6'd64,6'd66,6'd67,6'd69: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd62,6'd65,6'd68,6'd70,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd86: Enemy_img = 4'd6;
//6'd72,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd42,6'd46,6'd47,6'd52,6'd55,6'd58,6'd69,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd72,6'd73,6'd74,6'd75,6'd77,6'd86,6'd87: Enemy_img = 4'd6;
//6'd71,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd40,6'd41,6'd44,6'd45,6'd46,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd67: Enemy_img = 4'd14;
//6'd42,6'd47,6'd48,6'd51,6'd60,6'd65,6'd66,6'd68,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd70,6'd71,6'd72,6'd73,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd39,6'd74: Enemy_img = 4'd7;
//6'd40,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd53,6'd55,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd41,6'd42,6'd47,6'd51,6'd52,6'd64,6'd67,6'd80,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd69,6'd71,6'd72,6'd86,6'd89,6'd90,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd70,6'd73,6'd91: Enemy_img = 4'd7;
//6'd41,6'd43,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd57,6'd59,6'd61,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd44,6'd46,6'd52,6'd63,6'd78,6'd79,6'd83,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd72,6'd93,6'd94: Enemy_img = 4'd6;
//6'd39,6'd68,6'd69,6'd70,6'd71,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd41,6'd45,6'd51,6'd76,6'd79,6'd83,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd71,6'd94: Enemy_img = 4'd6;
//6'd39,6'd67,6'd68,6'd69,6'd70,6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd46,6'd50,6'd75,6'd76,6'd78,6'd82,6'd83,6'd86,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd93: Enemy_img = 4'd6;
//6'd39,6'd40,6'd69,6'd70,6'd92: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd48,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd67: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd74,6'd75,6'd77,6'd78,6'd83,6'd85,6'd86,6'd97,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38: Enemy_img = 4'd6;
//6'd39,6'd40,6'd69: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd45,6'd48,6'd68,6'd73,6'd74,6'd76,6'd77,6'd78,6'd82,6'd84,6'd85,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38: Enemy_img = 4'd6;
//6'd39,6'd40: Enemy_img = 4'd7;
//6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd44,6'd49,6'd66,6'd67,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd82,6'd83,6'd86,6'd87,6'd89,6'd93,6'd96,6'd98,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd2;
//6'd36,6'd37,6'd38: Enemy_img = 4'd6;
//6'd39,6'd40: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd67: Enemy_img = 4'd14;
//6'd44,6'd50,6'd65,6'd66,6'd70,6'd72,6'd73,6'd75,6'd76,6'd78,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd6;
//6'd38,6'd39: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd66: Enemy_img = 4'd14;
//6'd45,6'd51,6'd64,6'd65,6'd67,6'd68,6'd70,6'd71,6'd74,6'd77,6'd82,6'd83,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd95,6'd96,6'd98,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37: Enemy_img = 4'd6;
//6'd38,6'd39,6'd89,6'd90,6'd92,6'd93,6'd95: Enemy_img = 4'd7;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd65,6'd68: Enemy_img = 4'd14;
//6'd41,6'd42,6'd45,6'd46,6'd63,6'd64,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd82,6'd83,6'd87,6'd98,6'd99,6'd100,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd2;
//6'd34,6'd35,6'd36: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd7;
//6'd41,6'd42,6'd46,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd60,6'd67: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd47,6'd68,6'd69,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd101,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd62,6'd65: Enemy_img = 4'd2;
//6'd33,6'd34,6'd35,6'd36,6'd95,6'd97,6'd98,6'd99,6'd101: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd67,6'd68: Enemy_img = 4'd14;
//6'd44,6'd47,6'd48,6'd69,6'd75,6'd76,6'd77,6'd78,6'd103,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd2;
//6'd32,6'd33,6'd34,6'd35,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd101: Enemy_img = 4'd6;
//6'd36,6'd37,6'd38,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68: Enemy_img = 4'd14;
//6'd46,6'd47,6'd60,6'd61,6'd66,6'd69,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd2;
//6'd31,6'd32,6'd33,6'd34,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd6;
//6'd35,6'd36,6'd37,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd49,6'd51,6'd54,6'd55,6'd56,6'd63,6'd64,6'd66,6'd69: Enemy_img = 4'd14;
//6'd60,6'd61,6'd65,6'd67,6'd68,6'd70,6'd73,6'd74,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd2;
//6'd29,6'd30,6'd31,6'd32,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd53: Enemy_img = 4'd9;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd49,6'd50,6'd54,6'd55,6'd56,6'd68,6'd69: Enemy_img = 4'd14;
//6'd64,6'd65,6'd66,6'd67,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd28,6'd29,6'd30,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd52: Enemy_img = 4'd9;
//6'd42,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd65,6'd67,6'd69: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd57,6'd60,6'd63,6'd64,6'd66,6'd68,6'd70,6'd71,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd52,6'd53: Enemy_img = 4'd9;
//6'd41,6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd56,6'd58,6'd59,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70: Enemy_img = 4'd14;
//6'd23,6'd24,6'd25,6'd38,6'd39,6'd40,6'd42,6'd57,6'd60,6'd61,6'd62,6'd63,6'd69,6'd73,6'd74,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd53,6'd54: Enemy_img = 4'd10;
//6'd24,6'd25,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd38,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd55: Enemy_img = 4'd9;
//6'd54: Enemy_img = 4'd10;
//6'd25,6'd26,6'd27,6'd29,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//6'd24,6'd28,6'd30,6'd33,6'd62,6'd63,6'd65,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd55: Enemy_img = 4'd9;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd60,6'd61: Enemy_img = 4'd14;
//6'd33,6'd56,6'd58,6'd62,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd56: Enemy_img = 4'd9;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd14;
//6'd25,6'd52,6'd53,6'd57,6'd60,6'd61,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd56: Enemy_img = 4'd14;
//6'd51,6'd52,6'd57,6'd59,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd82,6'd83: Enemy_img = 4'd7;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd25,6'd26,6'd50,6'd51,6'd56,6'd57,6'd58,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd81,6'd82: Enemy_img = 4'd7;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd51,6'd52,6'd53,6'd54,6'd57: Enemy_img = 4'd14;
//6'd26,6'd27,6'd49,6'd50,6'd55,6'd56,6'd58,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd74,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd46,6'd84,6'd85: Enemy_img = 4'd6;
//6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd50,6'd51,6'd52,6'd56,6'd57: Enemy_img = 4'd14;
//6'd48,6'd49,6'd53,6'd54,6'd55,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd82: Enemy_img = 4'd7;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd51,6'd53,6'd54,6'd56,6'd57: Enemy_img = 4'd14;
//6'd27,6'd49,6'd50,6'd52,6'd55,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd47,6'd48,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd82: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd53,6'd55,6'd57: Enemy_img = 4'd14;
//6'd28,6'd50,6'd52,6'd54,6'd56,6'd58,6'd60,6'd61,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd76,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd47,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd57: Enemy_img = 4'd14;
//6'd54,6'd56,6'd60,6'd61,6'd62,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd47,6'd48,6'd83,6'd84: Enemy_img = 4'd6;
//6'd40,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Enemy_img = 4'd14;
//6'd28,6'd29,6'd49,6'd50,6'd58,6'd60,6'd61,6'd62,6'd63,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd46,6'd47,6'd83,6'd84: Enemy_img = 4'd6;
//6'd39,6'd40,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Enemy_img = 4'd14;
//6'd29,6'd30,6'd49,6'd50,6'd51,6'd60,6'd61,6'd62,6'd65,6'd66,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd83: Enemy_img = 4'd6;
//6'd38,6'd39,6'd43: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd52,6'd53,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd30,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd57,6'd58,6'd59,6'd60,6'd63,6'd65,6'd71,6'd73,6'd74,6'd77,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd83: Enemy_img = 4'd6;
//6'd37,6'd43,6'd44,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd7;
//6'd32,6'd33: Enemy_img = 4'd14;
//6'd30,6'd31,6'd46,6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd74,6'd76,6'd77,6'd79,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd39,6'd40,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd6;
//6'd37,6'd38,6'd41,6'd42,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd7;
//6'd31,6'd32: Enemy_img = 4'd14;
//6'd30,6'd44,6'd45,6'd48,6'd49,6'd51,6'd52,6'd54,6'd55,6'd56,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd39,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd30,6'd31,6'd43,6'd44,6'd45,6'd47,6'd53,6'd55,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd74,6'd77: Enemy_img = 4'd6;
//6'd36,6'd37,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd46,6'd47,6'd49,6'd51,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd6;
//6'd37,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd6;
//6'd56: Enemy_img = 4'd7;
//6'd39,6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58: Enemy_img = 4'd6;
//6'd56: Enemy_img = 4'd7;
//6'd43,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57: Enemy_img = 4'd6;
//6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55: Enemy_img = 4'd15;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd14;
//6'd83,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83,6'd84: Enemy_img = 4'd14;
//6'd81,6'd82,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd66,6'd80,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd13;
//6'd67,6'd68,6'd70,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd66,6'd78,6'd79,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd13;
//6'd67,6'd68,6'd70,6'd71,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd65,6'd66,6'd72,6'd76,6'd84,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd66,6'd67,6'd69,6'd70,6'd71,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd65,6'd72,6'd73,6'd75,6'd76,6'd77,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd66,6'd67,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd72,6'd73,6'd83,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd69,6'd70,6'd72,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd69,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd51,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73,6'd82,6'd83,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78,6'd79,6'd82: Enemy_img = 4'd6;
//6'd49,6'd52,6'd53,6'd58,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd59,6'd64,6'd67,6'd68,6'd71,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd82: Enemy_img = 4'd6;
//6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd68,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd51,6'd55,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd79,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd77,6'd78: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd91,6'd92: Enemy_img = 4'd14;
//6'd62,6'd63,6'd66,6'd67,6'd85,6'd86,6'd87,6'd88,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd79,6'd80: Enemy_img = 4'd6;
//6'd78,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd93: Enemy_img = 4'd13;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd65,6'd66,6'd69,6'd70,6'd74,6'd75,6'd76,6'd91,6'd92,6'd94: Enemy_img = 4'd14;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd67,6'd68,6'd71,6'd72,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd62,6'd79,6'd80: Enemy_img = 4'd6;
//6'd81,6'd82: Enemy_img = 4'd7;
//6'd93: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd70,6'd74,6'd75,6'd76,6'd77,6'd92,6'd94,6'd95: Enemy_img = 4'd14;
//6'd57,6'd58,6'd59,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd71,6'd72,6'd85,6'd87,6'd88,6'd89,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd60,6'd61,6'd62,6'd78,6'd79: Enemy_img = 4'd6;
//6'd51,6'd52,6'd67: Enemy_img = 4'd7;
//6'd92: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55,6'd56,6'd72,6'd74,6'd75,6'd76,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//6'd57,6'd58,6'd64,6'd68,6'd69,6'd70,6'd71,6'd73,6'd83,6'd84,6'd85,6'd89,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd59,6'd60,6'd61,6'd63,6'd78,6'd79: Enemy_img = 4'd6;
//6'd52,6'd62,6'd65,6'd66,6'd67: Enemy_img = 4'd7;
//6'd55,6'd56,6'd71,6'd72,6'd75,6'd76,6'd93,6'd94: Enemy_img = 4'd14;
//6'd57,6'd69,6'd70,6'd83,6'd84,6'd87,6'd88,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd63,6'd77,6'd78: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79: Enemy_img = 4'd7;
//6'd55,6'd94: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd70,6'd71,6'd72,6'd73,6'd75,6'd81,6'd83,6'd84,6'd85,6'd90,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd63,6'd64,6'd78: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd77: Enemy_img = 4'd7;
//6'd55,6'd56: Enemy_img = 4'd14;
//6'd57,6'd58,6'd59,6'd70,6'd71,6'd72,6'd73,6'd74,6'd80,6'd84,6'd89,6'd90,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd64,6'd69,6'd77,6'd78: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd60,6'd65,6'd66,6'd67,6'd68,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd56,6'd57: Enemy_img = 4'd14;
//6'd58,6'd59,6'd81,6'd85,6'd86,6'd87,6'd88,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd65,6'd72,6'd73,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd57: Enemy_img = 4'd14;
//6'd58,6'd59,6'd61,6'd62,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd78: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd76,6'd77,6'd79: Enemy_img = 4'd7;
//6'd58: Enemy_img = 4'd14;
//6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd83,6'd84,6'd86,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd64,6'd65,6'd72,6'd78,6'd79: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd58,6'd60,6'd61: Enemy_img = 4'd14;
//6'd57,6'd59,6'd62,6'd63,6'd68,6'd69,6'd89,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd78,6'd79: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd87: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd14;
//6'd63,6'd65,6'd66,6'd67,6'd68,6'd71,6'd91,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd79,6'd81: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66: Enemy_img = 4'd14;
//6'd64,6'd65,6'd67,6'd70,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd64: Enemy_img = 4'd14;
//6'd63,6'd65,6'd66,6'd67,6'd69,6'd70,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd82,6'd83,6'd91: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64: Enemy_img = 4'd14;
//6'd63,6'd65,6'd67,6'd68,6'd69,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd83,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd68: Enemy_img = 4'd14;
//6'd63,6'd64,6'd67,6'd69,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd71,6'd84,6'd86,6'd87,6'd88,6'd89,6'd91: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd72,6'd73,6'd74,6'd75,6'd76,6'd85,6'd90: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd61,6'd67: Enemy_img = 4'd14;
//6'd62,6'd63,6'd65,6'd66,6'd68,6'd69,6'd95,6'd96,6'd97,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd70,6'd71,6'd84,6'd85,6'd87,6'd92: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd72,6'd73,6'd74,6'd75,6'd76,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd58,6'd66,6'd67: Enemy_img = 4'd14;
//6'd57,6'd59,6'd60,6'd61,6'd64,6'd65,6'd68,6'd95,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd71,6'd74,6'd75,6'd84,6'd92: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd72,6'd73,6'd89,6'd90: Enemy_img = 4'd7;
//6'd64,6'd68: Enemy_img = 4'd14;
//6'd58,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd69,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd70,6'd71,6'd72,6'd74,6'd75: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd73,6'd89: Enemy_img = 4'd7;
//6'd62,6'd63,6'd65,6'd67: Enemy_img = 4'd14;
//6'd59,6'd60,6'd61,6'd64,6'd66,6'd68,6'd81,6'd95,6'd96,6'd99,6'd100,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd7;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd67: Enemy_img = 4'd14;
//6'd57,6'd58,6'd64,6'd65,6'd66,6'd68,6'd78,6'd82,6'd85,6'd86,6'd93,6'd94,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd104,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd71,6'd72,6'd73: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd70: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd62,6'd64: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd57,6'd61,6'd63,6'd65,6'd66,6'd67,6'd68,6'd76,6'd77,6'd82,6'd85,6'd90,6'd94,6'd95,6'd96,6'd99,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd69,6'd70,6'd71,6'd100,6'd102: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd72,6'd73,6'd95,6'd97,6'd98: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd54,6'd56,6'd61,6'd62,6'd63,6'd67,6'd78,6'd82,6'd84,6'd87,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd69,6'd70,6'd71,6'd99,6'd100: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd72,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd55,6'd56,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd60,6'd67,6'd75,6'd77,6'd78,6'd82,6'd86,6'd87,6'd88,6'd89,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd68,6'd69,6'd70,6'd71,6'd72,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd43,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd7;
//6'd50,6'd53,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd51,6'd54,6'd55,6'd58,6'd64,6'd65,6'd66,6'd75,6'd77,6'd78,6'd82,6'd83,6'd84,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68,6'd71,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd69,6'd70,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd7;
//6'd47,6'd49,6'd53,6'd54,6'd56,6'd58,6'd61,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd50,6'd51,6'd55,6'd57,6'd64,6'd74,6'd75,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd68,6'd69,6'd70,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd33,6'd34,6'd37,6'd39,6'd42,6'd45,6'd46,6'd47,6'd48,6'd51,6'd53,6'd54,6'd58,6'd61,6'd62,6'd64,6'd65: Enemy_img = 4'd14;
//6'd35,6'd36,6'd38,6'd40,6'd41,6'd43,6'd44,6'd49,6'd52,6'd55,6'd56,6'd57,6'd59,6'd60,6'd63,6'd74,6'd77,6'd78,6'd79,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd67,6'd69,6'd70,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd51,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd37,6'd43,6'd48,6'd50,6'd52,6'd53,6'd54,6'd74,6'd75,6'd76,6'd79,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd70,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd35,6'd44,6'd45,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd68: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd50,6'd51,6'd52,6'd72,6'd73,6'd74,6'd77,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd37,6'd38,6'd40,6'd41,6'd44,6'd45,6'd48,6'd49,6'd50,6'd52,6'd53,6'd55,6'd60,6'd62,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd39,6'd42,6'd43,6'd46,6'd51,6'd69,6'd74,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd39,6'd44,6'd46,6'd51,6'd52,6'd68,6'd69,6'd71,6'd72,6'd73,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd42,6'd46,6'd49,6'd50,6'd51,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd43,6'd47,6'd48,6'd52,6'd53,6'd68,6'd70,6'd72,6'd73,6'd74,6'd75,6'd77,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd68: Enemy_img = 4'd14;
//6'd42,6'd48,6'd52,6'd67,6'd69,6'd70,6'd71,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd2;
//6'd37,6'd38,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd68,6'd70: Enemy_img = 4'd14;
//6'd43,6'd47,6'd52,6'd67,6'd69,6'd71,6'd72,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64: Enemy_img = 4'd2;
//6'd37,6'd38,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd41,6'd42,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd68,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd43,6'd45,6'd46,6'd47,6'd51,6'd66,6'd67,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd2;
//6'd38,6'd39,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd40,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd41,6'd42,6'd44,6'd45,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd43,6'd46,6'd47,6'd48,6'd51,6'd73,6'd74,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67: Enemy_img = 4'd2;
//6'd38,6'd39,6'd40,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd69,6'd73: Enemy_img = 4'd14;
//6'd43,6'd48,6'd49,6'd50,6'd51,6'd70,6'd71,6'd72,6'd74,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd41,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd49,6'd50,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd43,6'd48,6'd51,6'd52,6'd53,6'd72,6'd75,6'd78,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd2;
//6'd39,6'd40,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd41,6'd42,6'd88,6'd89: Enemy_img = 4'd7;
//6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd57,6'd58,6'd59,6'd60,6'd64,6'd67,6'd68,6'd75: Enemy_img = 4'd14;
//6'd47,6'd48,6'd54,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd80,6'd81,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62: Enemy_img = 4'd2;
//6'd39,6'd40,6'd41,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd42,6'd43,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd47,6'd64,6'd69,6'd74,6'd75,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd65,6'd66: Enemy_img = 4'd2;
//6'd40,6'd41,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd42,6'd43,6'd88,6'd89: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd68,6'd73,6'd74,6'd78,6'd81,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64: Enemy_img = 4'd2;
//6'd40,6'd41,6'd42,6'd91,6'd92: Enemy_img = 4'd6;
//6'd43,6'd44,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd67,6'd69,6'd70: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd68,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd91,6'd92: Enemy_img = 4'd6;
//6'd43,6'd44,6'd89,6'd90: Enemy_img = 4'd7;
//6'd46,6'd48,6'd50,6'd51,6'd53,6'd54,6'd55,6'd57,6'd60,6'd61,6'd62,6'd64,6'd65,6'd69: Enemy_img = 4'd14;
//6'd47,6'd49,6'd52,6'd66,6'd67,6'd68,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd91,6'd92: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd90: Enemy_img = 4'd7;
//6'd58: Enemy_img = 4'd9;
//6'd46,6'd50,6'd51,6'd53,6'd54,6'd56,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd45,6'd47,6'd48,6'd49,6'd52,6'd63,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd92,6'd93: Enemy_img = 4'd6;
//6'd43,6'd44: Enemy_img = 4'd7;
//6'd58,6'd59: Enemy_img = 4'd9;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd56,6'd57,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd14;
//6'd52,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd91,6'd92: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44: Enemy_img = 4'd7;
//6'd59,6'd60,6'd62: Enemy_img = 4'd9;
//6'd61: Enemy_img = 4'd10;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd67,6'd68,6'd72,6'd73,6'd74,6'd75,6'd78,6'd79,6'd80,6'd81,6'd85,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd92,6'd93: Enemy_img = 4'd6;
//6'd43,6'd44: Enemy_img = 4'd7;
//6'd63: Enemy_img = 4'd9;
//6'd60,6'd61,6'd62: Enemy_img = 4'd10;
//6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd64,6'd65,6'd67,6'd73,6'd74,6'd75,6'd77,6'd81,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd6;
//6'd43,6'd44: Enemy_img = 4'd7;
//6'd62,6'd63: Enemy_img = 4'd9;
//6'd46,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd14;
//6'd66,6'd67,6'd70,6'd71,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd93: Enemy_img = 4'd6;
//6'd42,6'd43: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd64: Enemy_img = 4'd14;
//6'd48,6'd61,6'd65,6'd66,6'd69,6'd70,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44: Enemy_img = 4'd7;
//6'd48,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd66: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd60,6'd65,6'd69,6'd70,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd85,6'd87,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd7;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd65,6'd66: Enemy_img = 4'd14;
//6'd46,6'd60,6'd64,6'd70,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd84,6'd87,6'd88,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd65,6'd66: Enemy_img = 4'd14;
//6'd59,6'd63,6'd64,6'd67,6'd69,6'd70,6'd71,6'd75,6'd76,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd67: Enemy_img = 4'd14;
//6'd59,6'd62,6'd64,6'd65,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd82,6'd83,6'd85,6'd87,6'd93,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd86,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd81,6'd83,6'd84: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67: Enemy_img = 4'd14;
//6'd59,6'd62,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd37,6'd38,6'd40,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd42,6'd43,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd71,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd56,6'd57,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd41,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd34,6'd36,6'd38,6'd39,6'd40,6'd42,6'd70,6'd71,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd58,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd56,6'd57,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd37,6'd67,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd58,6'd59,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd56,6'd57,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd33,6'd60,6'd61,6'd62,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd58,6'd59,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd51: Enemy_img = 4'd14;
//6'd34,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd58,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd72,6'd73: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51: Enemy_img = 4'd14;
//6'd34,6'd35,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd67,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd58,6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd56,6'd57,6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd52,6'd54,6'd55,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd52,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd14;
//6'd38,6'd59,6'd60,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd51,6'd52,6'd57,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd59,6'd60,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd73,6'd74,6'd75: Enemy_img = 4'd6;
//6'd51,6'd52,6'd55,6'd56,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd58,6'd65,6'd66,6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd73,6'd74: Enemy_img = 4'd6;
//6'd50,6'd55,6'd56,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd41,6'd42,6'd58,6'd59,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd74: Enemy_img = 4'd6;
//6'd55,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd58,6'd59,6'd61,6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd53,6'd54,6'd73: Enemy_img = 4'd6;
//6'd52,6'd55,6'd71,6'd72: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd43,6'd44,6'd57,6'd58,6'd60,6'd64,6'd65,6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd53,6'd54,6'd55,6'd74: Enemy_img = 4'd6;
//6'd51,6'd52,6'd72,6'd73: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd57,6'd58,6'd60,6'd61,6'd62,6'd64,6'd65,6'd67,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd53,6'd54,6'd74: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52: Enemy_img = 4'd7;
//6'd47: Enemy_img = 4'd14;
//6'd45,6'd46,6'd56,6'd57,6'd60,6'd61,6'd62,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd73: Enemy_img = 4'd6;
//6'd53: Enemy_img = 4'd7;
//6'd45,6'd46,6'd56,6'd57,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53: Enemy_img = 4'd6;
//6'd46,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd62,6'd65,6'd67,6'd68,6'd70,6'd71,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd14;
//6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd14;
//6'd66,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67: Enemy_img = 4'd14;
//6'd65,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd64,6'd68,6'd69,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd64,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd63,6'd68,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66: Enemy_img = 4'd14;
//6'd62,6'd67,6'd68,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd61,6'd68,6'd69,6'd70,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd61,6'd62,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd80: Enemy_img = 4'd13;
//6'd52,6'd53,6'd55,6'd56,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd14;
//6'd51,6'd57,6'd58,6'd60,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd77,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd80: Enemy_img = 4'd13;
//6'd52,6'd53,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd78,6'd79,6'd81,6'd82: Enemy_img = 4'd14;
//6'd51,6'd57,6'd59,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd69: Enemy_img = 4'd6;
//6'd54,6'd80: Enemy_img = 4'd13;
//6'd52,6'd53,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd81,6'd82: Enemy_img = 4'd14;
//6'd51,6'd58,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd6;
//6'd67,6'd68: Enemy_img = 4'd7;
//6'd54: Enemy_img = 4'd13;
//6'd52,6'd53,6'd60,6'd61,6'd62,6'd63,6'd81,6'd82: Enemy_img = 4'd14;
//6'd51,6'd56,6'd58,6'd59,6'd75,6'd76,6'd77,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd64,6'd65,6'd70,6'd71: Enemy_img = 4'd7;
//6'd52,6'd53,6'd59,6'd60,6'd61,6'd62,6'd82: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd73,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd7;
//6'd56,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd54,6'd55,6'd57,6'd72,6'd73,6'd75,6'd76,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd66,6'd69: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd58,6'd71,6'd72,6'd73,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd6;
//6'd67: Enemy_img = 4'd7;
//6'd54,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd72,6'd73,6'd74,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd55,6'd60,6'd70,6'd72,6'd73,6'd76,6'd77,6'd78,6'd80,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd6;
//6'd68: Enemy_img = 4'd7;
//6'd50,6'd51,6'd56,6'd58,6'd59,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd52,6'd53,6'd54,6'd55,6'd57,6'd60,6'd61,6'd70,6'd75,6'd76,6'd77,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd59,6'd61,6'd64,6'd65: Enemy_img = 4'd14;
//6'd45,6'd46,6'd47,6'd52,6'd56,6'd57,6'd58,6'd60,6'd62,6'd70,6'd71,6'd74,6'd75,6'd76,6'd80,6'd82,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd6;
//6'd67: Enemy_img = 4'd7;
//6'd46,6'd48,6'd49,6'd50,6'd54,6'd61,6'd62: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd47,6'd51,6'd52,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd63,6'd65,6'd73,6'd74,6'd75,6'd85,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd57,6'd66,6'd69,6'd78: Enemy_img = 4'd7;
//6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50,6'd51,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd87,6'd88,6'd89,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd66,6'd69,6'd83: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd65,6'd67,6'd68,6'd70,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd40,6'd44,6'd48,6'd49,6'd50,6'd54,6'd60,6'd61,6'd62,6'd63,6'd87,6'd88,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd65,6'd66,6'd69,6'd70,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd64,6'd67,6'd68,6'd71,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd39,6'd40,6'd48,6'd49,6'd88,6'd90,6'd91,6'd92,6'd93,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd53,6'd54,6'd60,6'd61,6'd62,6'd64,6'd65,6'd70,6'd71,6'd73,6'd74,6'd75,6'd81,6'd82,6'd84,6'd85: Enemy_img = 4'd6;
//6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd63,6'd66,6'd67,6'd68,6'd69,6'd72,6'd76,6'd77,6'd78,6'd79,6'd80,6'd83: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd47,6'd48,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd50,6'd54,6'd55,6'd59,6'd60,6'd62,6'd63,6'd64,6'd71,6'd72,6'd73,6'd75,6'd76,6'd80,6'd81,6'd85,6'd96: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd56,6'd57,6'd58,6'd61,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd77,6'd78,6'd79,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd14;
//6'd47,6'd48,6'd89,6'd90,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd55,6'd56,6'd58,6'd59,6'd76,6'd77,6'd79,6'd80,6'd94,6'd95: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd57,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd78,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd48,6'd49,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd56,6'd57,6'd58,6'd77,6'd78,6'd79,6'd94,6'd95: Enemy_img = 4'd6;
//6'd42,6'd43,6'd52,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd83,6'd92,6'd93: Enemy_img = 4'd7;
//6'd46: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd50,6'd54,6'd60,6'd61,6'd63,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd57,6'd78,6'd93,6'd94: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd47,6'd48,6'd49: Enemy_img = 4'd14;
//6'd50,6'd51,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd48,6'd49,6'd54: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd62,6'd63,6'd81,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd92,6'd93: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd49,6'd51,6'd53,6'd54,6'd55,6'd59: Enemy_img = 4'd14;
//6'd50,6'd52,6'd56,6'd57,6'd58,6'd60,6'd62,6'd63,6'd76,6'd80,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd65,6'd70,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd66,6'd67,6'd68,6'd69,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58: Enemy_img = 4'd14;
//6'd50,6'd57,6'd59,6'd61,6'd62,6'd63,6'd77,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd65,6'd66,6'd69,6'd70,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd67,6'd68,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd62: Enemy_img = 4'd14;
//6'd57,6'd59,6'd61,6'd63,6'd73,6'd77,6'd78,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd65,6'd66,6'd69,6'd70,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd67,6'd68,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd62: Enemy_img = 4'd14;
//6'd57,6'd58,6'd60,6'd61,6'd63,6'd73,6'd78,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd66,6'd67,6'd68,6'd69,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd58,6'd60,6'd64,6'd72,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd66,6'd67,6'd68,6'd69,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd63: Enemy_img = 4'd14;
//6'd57,6'd59,6'd60,6'd61,6'd62,6'd64,6'd74,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd67,6'd68,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd66,6'd69,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd60,6'd61,6'd63: Enemy_img = 4'd14;
//6'd56,6'd58,6'd59,6'd62,6'd64,6'd72,6'd74,6'd75,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd67,6'd68,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd66,6'd69,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd53,6'd54,6'd59,6'd63: Enemy_img = 4'd14;
//6'd55,6'd57,6'd58,6'd60,6'd61,6'd62,6'd64,6'd72,6'd74,6'd75,6'd76,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd66,6'd67,6'd68,6'd69,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd58,6'd59,6'd61: Enemy_img = 4'd14;
//6'd53,6'd54,6'd56,6'd57,6'd60,6'd62,6'd63,6'd64,6'd72,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd66,6'd67,6'd68,6'd69,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd55,6'd56,6'd60,6'd64,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd66,6'd69,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd67,6'd68,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd56,6'd57,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd54,6'd55,6'd58,6'd59,6'd60,6'd64,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd66,6'd69,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd67,6'd68,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//6'd54,6'd58,6'd62,6'd63,6'd64,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd66,6'd67,6'd68,6'd69,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd56,6'd57,6'd59,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd52,6'd58,6'd62,6'd71,6'd72,6'd73,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd66,6'd69,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd61,6'd63,6'd64: Enemy_img = 4'd14;
//6'd51,6'd52,6'd54,6'd55,6'd62,6'd75,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd60,6'd61,6'd63,6'd64,6'd67: Enemy_img = 4'd14;
//6'd50,6'd51,6'd56,6'd57,6'd62,6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd55,6'd57,6'd62,6'd63,6'd66,6'd67: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd53,6'd54,6'd56,6'd58,6'd59,6'd68,6'd69,6'd72,6'd73,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd69: Enemy_img = 4'd14;
//6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd68,6'd70,6'd71,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd49,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd71: Enemy_img = 4'd14;
//6'd47,6'd48,6'd50,6'd54,6'd68,6'd70,6'd72,6'd73,6'd78,6'd79,6'd80,6'd82,6'd83,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd94,6'd95: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd48,6'd51,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd46,6'd47,6'd49,6'd52,6'd53,6'd54,6'd68,6'd70,6'd74,6'd75,6'd80,6'd82,6'd83,6'd84,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd42,6'd93: Enemy_img = 4'd7;
//6'd47,6'd48,6'd51,6'd53,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd69,6'd72,6'd73,6'd75: Enemy_img = 4'd14;
//6'd45,6'd46,6'd49,6'd52,6'd68,6'd74,6'd76,6'd77,6'd82,6'd83,6'd84,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd70: Enemy_img = 4'd2;
//6'd39,6'd40,6'd95,6'd96: Enemy_img = 4'd6;
//6'd46,6'd47,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd67,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd48,6'd50,6'd51,6'd52,6'd68,6'd72,6'd73,6'd74,6'd78,6'd79,6'd84,6'd85,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd69: Enemy_img = 4'd2;
//6'd38,6'd39,6'd96,6'd97: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd50,6'd51,6'd53,6'd54,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd48,6'd52,6'd74,6'd75,6'd76,6'd77,6'd78,6'd81,6'd82,6'd84,6'd85,6'd88,6'd89,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd2;
//6'd37,6'd98: Enemy_img = 4'd6;
//6'd42,6'd43,6'd45,6'd46,6'd49,6'd50,6'd51,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd70,6'd71,6'd75,6'd76: Enemy_img = 4'd14;
//6'd40,6'd41,6'd44,6'd47,6'd52,6'd53,6'd54,6'd72,6'd73,6'd74,6'd77,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd38,6'd39,6'd44,6'd47,6'd54,6'd72,6'd76,6'd79,6'd80,6'd81,6'd82,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd45,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd73,6'd74: Enemy_img = 4'd14;
//6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd46,6'd48,6'd49,6'd50,6'd54,6'd68,6'd69,6'd72,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd70: Enemy_img = 4'd2;
//6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd67,6'd73,6'd74: Enemy_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd46,6'd50,6'd54,6'd68,6'd72,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd90,6'd91,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd69: Enemy_img = 4'd2;
//6'd36,6'd37,6'd39,6'd40,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd71,6'd73: Enemy_img = 4'd14;
//6'd38,6'd41,6'd45,6'd50,6'd54,6'd72,6'd74,6'd77,6'd78,6'd79,6'd80,6'd88,6'd91,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd2;
//6'd39,6'd40,6'd47,6'd48,6'd49,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd50,6'd54,6'd70,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd93,6'd94,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd97: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd41,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd74,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd95,6'd96: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73: Enemy_img = 4'd14;
//6'd46,6'd52,6'd68,6'd74,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd45,6'd46,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd14;
//6'd47,6'd52,6'd73,6'd76,6'd77,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd44,6'd91: Enemy_img = 4'd7;
//6'd64: Enemy_img = 4'd9;
//6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62: Enemy_img = 4'd14;
//6'd47,6'd52,6'd71,6'd73,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd45,6'd46,6'd89,6'd90: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd9;
//6'd67: Enemy_img = 4'd10;
//6'd50,6'd51,6'd59,6'd60,6'd62: Enemy_img = 4'd14;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd70,6'd71,6'd73,6'd76,6'd77,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd65,6'd69,6'd70: Enemy_img = 4'd9;
//6'd66,6'd67,6'd68: Enemy_img = 4'd10;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63: Enemy_img = 4'd14;
//6'd55,6'd58,6'd72,6'd73,6'd76,6'd77,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd89,6'd90,6'd91: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd59,6'd61,6'd62,6'd63,6'd64,6'd71,6'd73: Enemy_img = 4'd14;
//6'd55,6'd58,6'd72,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd52,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd73,6'd74: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd68,6'd69,6'd72,6'd75,6'd78,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd49,6'd50,6'd85,6'd86: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75: Enemy_img = 4'd14;
//6'd52,6'd68,6'd72,6'd76,6'd79,6'd80,6'd81,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd76: Enemy_img = 4'd14;
//6'd68,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd50,6'd51,6'd84,6'd85: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd68,6'd71,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd68,6'd71,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd51,6'd52,6'd83,6'd84: Enemy_img = 4'd7;
//6'd54,6'd55,6'd59,6'd60,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd68,6'd71,6'd72,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd51,6'd52,6'd83,6'd84: Enemy_img = 4'd7;
//6'd54,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67: Enemy_img = 4'd14;
//6'd55,6'd56,6'd68,6'd69,6'd70,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd55,6'd73,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd66,6'd67,6'd68,6'd69,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd14;
//6'd55,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd65,6'd66,6'd69,6'd70,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd67,6'd68,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd65,6'd66,6'd69,6'd70,6'd86,6'd87: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd67,6'd68,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd72,6'd73,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd65,6'd70,6'd86,6'd87: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd66,6'd67,6'd68,6'd69,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd72,6'd73,6'd75,6'd76,6'd77,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd65,6'd70,6'd87: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd66,6'd67,6'd68,6'd69,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd54,6'd72,6'd73,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd65,6'd66,6'd69,6'd70,6'd87,6'd88: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd67,6'd68,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd54,6'd55,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd53,6'd72,6'd73,6'd75,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd65,6'd66,6'd69,6'd70,6'd88: Enemy_img = 4'd6;
//6'd48,6'd49,6'd67,6'd68,6'd86,6'd87: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63: Enemy_img = 4'd14;
//6'd52,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd66,6'd67,6'd68,6'd69,6'd88: Enemy_img = 4'd6;
//6'd65,6'd70: Enemy_img = 4'd7;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd14;
//6'd50,6'd51,6'd75,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd65,6'd70: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd48,6'd49,6'd72,6'd73,6'd75,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd7;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd46,6'd47,6'd72,6'd73,6'd75,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67,6'd68: Enemy_img = 4'd6;
//6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd7;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd44,6'd45,6'd72,6'd73,6'd75,6'd76,6'd77,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd65,6'd70: Enemy_img = 4'd7;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd46,6'd47,6'd72,6'd73,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd6;
//6'd65,6'd70: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd48,6'd49,6'd72,6'd73,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd6;
//6'd67,6'd68: Enemy_img = 4'd7;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd72,6'd73,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd69,6'd70: Enemy_img = 4'd6;
//6'd67,6'd68: Enemy_img = 4'd7;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd72,6'd73,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd70: Enemy_img = 4'd6;
//6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd7;
//6'd59,6'd60,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd56,6'd57,6'd58,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd70: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd59,6'd60,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd14;
//6'd61,6'd62,6'd72,6'd73,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63: Enemy_img = 4'd15;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd14;
//6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52: Enemy_img = 4'd14;
//6'd51,6'd53,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd14;
//6'd53,6'd54,6'd55,6'd56,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd68,6'd69: Enemy_img = 4'd14;
//6'd54,6'd57,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd67: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd65,6'd66,6'd68,6'd69: Enemy_img = 4'd14;
//6'd50,6'd54,6'd56,6'd59,6'd60,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd68: Enemy_img = 4'd13;
//6'd51,6'd52,6'd53,6'd65,6'd66,6'd67,6'd69,6'd70: Enemy_img = 4'd14;
//6'd50,6'd54,6'd55,6'd57,6'd59,6'd64,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd69,6'd70: Enemy_img = 4'd14;
//6'd50,6'd54,6'd55,6'd56,6'd60,6'd61,6'd62,6'd63,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd49,6'd56,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd49,6'd50,6'd56,6'd59,6'd60,6'd68,6'd69,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd58,6'd59: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd14;
//6'd49,6'd62,6'd64,6'd65,6'd67,6'd68,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd82,6'd84,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd58: Enemy_img = 4'd6;
//6'd56,6'd57,6'd59,6'd60: Enemy_img = 4'd7;
//6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd14;
//6'd48,6'd61,6'd62,6'd63,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd88: Enemy_img = 4'd6;
//6'd59,6'd60: Enemy_img = 4'd7;
//6'd45,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd70,6'd71,6'd73,6'd76,6'd78,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd87: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd59: Enemy_img = 4'd7;
//6'd43: Enemy_img = 4'd13;
//6'd44,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd46,6'd62,6'd63,6'd67,6'd68,6'd71,6'd78,6'd79,6'd80,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd75,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd55,6'd56: Enemy_img = 4'd7;
//6'd43: Enemy_img = 4'd13;
//6'd41,6'd42,6'd44,6'd45,6'd50,6'd51,6'd52: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd63,6'd66,6'd67,6'd82,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd75,6'd76,6'd77,6'd87: Enemy_img = 4'd6;
//6'd58,6'd70,6'd85,6'd86: Enemy_img = 4'd7;
//6'd44: Enemy_img = 4'd13;
//6'd41,6'd42,6'd43,6'd45,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd56: Enemy_img = 4'd14;
//6'd40,6'd46,6'd48,6'd61,6'd65,6'd66,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd74,6'd76,6'd77,6'd78,6'd86,6'd87: Enemy_img = 4'd6;
//6'd59,6'd70,6'd71,6'd72,6'd75,6'd85: Enemy_img = 4'd7;
//6'd44: Enemy_img = 4'd13;
//6'd42,6'd43,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd41,6'd46,6'd47,6'd61,6'd62,6'd65,6'd66,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd74,6'd86,6'd87: Enemy_img = 4'd6;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd42,6'd43,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd41,6'd45,6'd46,6'd48,6'd49,6'd80,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd73,6'd74,6'd86,6'd87: Enemy_img = 4'd6;
//6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd43,6'd47,6'd48,6'd53,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd45,6'd46,6'd49,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd68,6'd73,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd59,6'd61,6'd62,6'd63,6'd69,6'd70,6'd71,6'd72,6'd77,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd46,6'd49,6'd50,6'd51,6'd56: Enemy_img = 4'd14;
//6'd44,6'd45,6'd47,6'd48,6'd52,6'd53,6'd57,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd64,6'd65,6'd72,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd46,6'd48,6'd49,6'd50,6'd51,6'd53: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd47,6'd52,6'd54,6'd55,6'd57,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd58,6'd60,6'd61,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd45,6'd46,6'd48,6'd51,6'd54: Enemy_img = 4'd14;
//6'd43,6'd44,6'd47,6'd49,6'd50,6'd52,6'd53,6'd55,6'd56,6'd57,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd65,6'd72,6'd73,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd47,6'd48: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd50,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd43,6'd44,6'd46,6'd47: Enemy_img = 4'd14;
//6'd41,6'd42,6'd45,6'd48,6'd49,6'd52,6'd53,6'd54,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd58,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd82,6'd83,6'd84: Enemy_img = 4'd7;
//6'd43,6'd44,6'd47: Enemy_img = 4'd14;
//6'd40,6'd41,6'd42,6'd45,6'd46,6'd48,6'd71,6'd75,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd40,6'd44,6'd45,6'd47,6'd48,6'd73,6'd74,6'd76,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd54,6'd55,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd40,6'd42,6'd43: Enemy_img = 4'd14;
//6'd38,6'd39,6'd41,6'd44,6'd45,6'd73,6'd74,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49,6'd54,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd38,6'd39,6'd43,6'd44,6'd56,6'd58,6'd69,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd48,6'd49,6'd50,6'd51,6'd53,6'd66,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd47,6'd52,6'd61,6'd62,6'd63,6'd64,6'd65,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd42,6'd43,6'd44,6'd55,6'd56,6'd57,6'd59,6'd70,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd50,6'd52,6'd53,6'd66,6'd67,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd61,6'd62,6'd63,6'd64,6'd65,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd38,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd36,6'd37,6'd39,6'd43,6'd55,6'd56,6'd58,6'd59,6'd70,6'd71,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd53,6'd62,6'd63,6'd66,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd47,6'd48,6'd64,6'd65,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd34,6'd35,6'd42,6'd43,6'd50,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd69,6'd71,6'd72,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd65,6'd66,6'd67,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd48,6'd64,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd56: Enemy_img = 4'd14;
//6'd35,6'd43,6'd44,6'd45,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd58,6'd59,6'd60,6'd70,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd51,6'd52,6'd55,6'd59: Enemy_img = 4'd14;
//6'd34,6'd35,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd53,6'd54,6'd56,6'd58,6'd60,6'd62,6'd70,6'd72,6'd73,6'd74,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd67,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd36,6'd38,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd50,6'd51,6'd52,6'd53,6'd55,6'd60,6'd61: Enemy_img = 4'd14;
//6'd43,6'd47,6'd48,6'd49,6'd54,6'd56,6'd58,6'd59,6'd62,6'd71,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd35,6'd37,6'd66,6'd67,6'd68,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd39,6'd40,6'd42,6'd64,6'd65,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd61: Enemy_img = 4'd14;
//6'd47,6'd49,6'd55,6'd56,6'd58,6'd60,6'd62,6'd71,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd66,6'd67,6'd68,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd65,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd60,6'd62: Enemy_img = 4'd14;
//6'd48,6'd56,6'd58,6'd59,6'd61,6'd63,6'd71,6'd72,6'd73,6'd77,6'd78,6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd39,6'd40,6'd65,6'd66,6'd67,6'd68,6'd69,6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd94: Enemy_img = 4'd7;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd62: Enemy_img = 4'd14;
//6'd56,6'd58,6'd61,6'd63,6'd72,6'd73,6'd75,6'd77,6'd80,6'd81,6'd84,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd66,6'd69: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd67,6'd68: Enemy_img = 4'd7;
//6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd63: Enemy_img = 4'd14;
//6'd57,6'd59,6'd60,6'd61,6'd62,6'd64,6'd71,6'd72,6'd73,6'd75,6'd76,6'd79,6'd80,6'd81,6'd83,6'd84,6'd88,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd66: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd67,6'd68,6'd69: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd60,6'd64,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd89,6'd90,6'd91,6'd93,6'd95,6'd98,6'd100,6'd103,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd67,6'd68,6'd70: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd61,6'd62,6'd63: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd60,6'd64,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd67: Enemy_img = 4'd7;
//6'd53,6'd57,6'd58,6'd61,6'd62,6'd64,6'd65: Enemy_img = 4'd14;
//6'd54,6'd56,6'd59,6'd60,6'd63,6'd69,6'd73,6'd74,6'd84,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd96,6'd97,6'd100,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd7;
//6'd57,6'd58,6'd60,6'd61,6'd62,6'd64,6'd65,6'd68,6'd69: Enemy_img = 4'd14;
//6'd53,6'd55,6'd56,6'd59,6'd63,6'd70,6'd71,6'd72,6'd73,6'd75,6'd77,6'd85,6'd87,6'd88,6'd89,6'd92,6'd93,6'd94,6'd95,6'd98,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd101: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd7;
//6'd57,6'd58,6'd60,6'd61,6'd62,6'd65,6'd66,6'd68,6'd69,6'd71,6'd73,6'd75,6'd78,6'd80: Enemy_img = 4'd14;
//6'd55,6'd56,6'd59,6'd63,6'd64,6'd70,6'd72,6'd74,6'd76,6'd77,6'd79,6'd81,6'd82,6'd84,6'd85,6'd87,6'd94,6'd95,6'd97,6'd98,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd101: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Enemy_img = 4'd7;
//6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd71,6'd74,6'd75,6'd76,6'd78,6'd79: Enemy_img = 4'd14;
//6'd55,6'd64,6'd70,6'd72,6'd73,6'd77,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd95,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd100: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd7;
//6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd54,6'd57,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd2;
//6'd44,6'd45,6'd46,6'd99,6'd100: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Enemy_img = 4'd7;
//6'd57,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd54,6'd56,6'd58,6'd59,6'd60,6'd61,6'd71,6'd75,6'd78,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd99,6'd100: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd58,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd53,6'd54,6'd59,6'd72,6'd76,6'd77,6'd80,6'd82,6'd83,6'd84,6'd85,6'd89,6'd90,6'd91,6'd92,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd98,6'd99: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd97: Enemy_img = 4'd7;
//6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd76,6'd80,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd71,6'd72: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd48,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51: Enemy_img = 4'd7;
//6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd53,6'd54,6'd57,6'd77,6'd80,6'd82,6'd83,6'd84,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd96: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd78: Enemy_img = 4'd14;
//6'd52,6'd53,6'd58,6'd74,6'd77,6'd79,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd97,6'd98: Enemy_img = 4'd6;
//6'd48,6'd49,6'd95,6'd96: Enemy_img = 4'd7;
//6'd53,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd77: Enemy_img = 4'd14;
//6'd52,6'd54,6'd56,6'd57,6'd73,6'd78,6'd79,6'd80,6'd83,6'd85,6'd86,6'd88,6'd89,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd94,6'd95: Enemy_img = 4'd7;
//6'd55,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd73,6'd79: Enemy_img = 4'd14;
//6'd51,6'd52,6'd53,6'd56,6'd77,6'd78,6'd80,6'd86,6'd87,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd74: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd96,6'd97: Enemy_img = 4'd6;
//6'd48,6'd49,6'd94,6'd95: Enemy_img = 4'd7;
//6'd52,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd51,6'd53,6'd54,6'd56,6'd57,6'd76,6'd81,6'd83,6'd84,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd2;
//6'd45,6'd46,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd93,6'd94: Enemy_img = 4'd7;
//6'd52,6'd53,6'd56,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd51,6'd55,6'd57,6'd59,6'd80,6'd83,6'd84,6'd86,6'd87,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd47,6'd48,6'd93,6'd94: Enemy_img = 4'd7;
//6'd51,6'd52,6'd55,6'd56,6'd57,6'd59,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77: Enemy_img = 4'd14;
//6'd50,6'd53,6'd58,6'd60,6'd75,6'd80,6'd84,6'd85,6'd88,6'd89,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd96,6'd97: Enemy_img = 4'd6;
//6'd47,6'd93,6'd94,6'd95: Enemy_img = 4'd7;
//6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd49,6'd50,6'd60,6'd79,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd93,6'd94: Enemy_img = 4'd7;
//6'd51,6'd52,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74: Enemy_img = 4'd14;
//6'd49,6'd50,6'd53,6'd61,6'd78,6'd79,6'd80,6'd81,6'd85,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd96,6'd97: Enemy_img = 4'd6;
//6'd93,6'd94,6'd95: Enemy_img = 4'd7;
//6'd76,6'd77,6'd78: Enemy_img = 4'd9;
//6'd75: Enemy_img = 4'd10;
//6'd49,6'd51,6'd52,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd66,6'd69,6'd70,6'd82,6'd83: Enemy_img = 4'd14;
//6'd47,6'd48,6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61,6'd65,6'd80,6'd81,6'd84,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd93,6'd94: Enemy_img = 4'd7;
//6'd72,6'd73,6'd74: Enemy_img = 4'd9;
//6'd75,6'd76,6'd77: Enemy_img = 4'd10;
//6'd48,6'd49,6'd50,6'd52,6'd55,6'd56,6'd58,6'd59,6'd60,6'd65,6'd66,6'd67,6'd68,6'd70,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd47,6'd51,6'd53,6'd57,6'd61,6'd62,6'd63,6'd64,6'd81,6'd85,6'd86,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd93,6'd94: Enemy_img = 4'd7;
//6'd74: Enemy_img = 4'd9;
//6'd75: Enemy_img = 4'd10;
//6'd47,6'd48,6'd49,6'd52,6'd55,6'd56,6'd59,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd71,6'd79,6'd80,6'd82,6'd83: Enemy_img = 4'd14;
//6'd50,6'd51,6'd53,6'd57,6'd58,6'd60,6'd61,6'd62,6'd78,6'd81,6'd84,6'd85,6'd86,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd94,6'd95: Enemy_img = 4'd7;
//6'd47,6'd50,6'd51,6'd55,6'd56,6'd57,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd76,6'd79,6'd80,6'd84: Enemy_img = 4'd14;
//6'd45,6'd46,6'd48,6'd49,6'd52,6'd53,6'd58,6'd59,6'd60,6'd77,6'd78,6'd81,6'd82,6'd83,6'd85,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd93,6'd94,6'd95: Enemy_img = 4'd7;
//6'd45,6'd46,6'd50,6'd51,6'd52,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd82,6'd83: Enemy_img = 4'd14;
//6'd47,6'd48,6'd49,6'd53,6'd56,6'd57,6'd60,6'd61,6'd66,6'd67,6'd78,6'd81,6'd84,6'd88,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd98,6'd99: Enemy_img = 4'd6;
//6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd7;
//6'd45,6'd48,6'd53,6'd57,6'd58,6'd59,6'd60,6'd62,6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd83: Enemy_img = 4'd14;
//6'd44,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52,6'd54,6'd61,6'd63,6'd64,6'd65,6'd67,6'd78,6'd81,6'd82,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd98,6'd99: Enemy_img = 4'd6;
//6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd60,6'd63,6'd64,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd46,6'd49,6'd55,6'd56,6'd61,6'd62,6'd65,6'd68,6'd79,6'd82,6'd83,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd100,6'd101: Enemy_img = 4'd6;
//6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd7;
//6'd42,6'd44,6'd52,6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81: Enemy_img = 4'd14;
//6'd50,6'd56,6'd65,6'd79,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd51,6'd101: Enemy_img = 4'd6;
//6'd53,6'd54,6'd56,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd64,6'd65,6'd79,6'd80,6'd81,6'd85,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd102: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd97,6'd99,6'd100: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd80,6'd81,6'd83: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72: Enemy_img = 4'd14;
//6'd63,6'd85,6'd86,6'd88,6'd89,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd79,6'd82,6'd83: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd80,6'd81: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd70,6'd85,6'd86,6'd92,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd78,6'd79,6'd82,6'd83: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63,6'd80,6'd81: Enemy_img = 4'd7;
//6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd68,6'd69,6'd85,6'd86,6'd87,6'd89,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61,6'd78,6'd79,6'd84: Enemy_img = 4'd6;
//6'd62,6'd63,6'd64,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd7;
//6'd66,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd86,6'd87,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60,6'd61,6'd62,6'd63,6'd79,6'd83,6'd84: Enemy_img = 4'd6;
//6'd64,6'd65,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd68,6'd86,6'd87,6'd90,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd79,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd68,6'd90,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd80,6'd81,6'd84: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66,6'd67,6'd82,6'd83,6'd85: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd14;
//6'd87,6'd88,6'd90,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd65,6'd66,6'd67,6'd85: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd87,6'd88,6'd89,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd65,6'd66,6'd67,6'd80,6'd85,6'd86: Enemy_img = 4'd7;
//6'd73,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd88,6'd89,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd83,6'd84: Enemy_img = 4'd6;
//6'd65,6'd66,6'd67,6'd68,6'd81,6'd82,6'd85,6'd86: Enemy_img = 4'd7;
//6'd70,6'd71,6'd72,6'd74,6'd76,6'd77,6'd79: Enemy_img = 4'd14;
//6'd69,6'd88,6'd89,6'd92,6'd93,6'd94,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd65,6'd66,6'd67,6'd81,6'd82,6'd87: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd89,6'd90,6'd92,6'd93,6'd94,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66,6'd67,6'd82: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd14;
//6'd89,6'd90,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd6;
//6'd65,6'd66,6'd82,6'd85: Enemy_img = 4'd7;
//6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd68,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd82,6'd83,6'd84,6'd87,6'd88: Enemy_img = 4'd6;
//6'd64,6'd65,6'd85,6'd86: Enemy_img = 4'd7;
//6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd67,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd83,6'd84,6'd88: Enemy_img = 4'd6;
//6'd85,6'd86,6'd87: Enemy_img = 4'd7;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd83: Enemy_img = 4'd6;
//6'd84: Enemy_img = 4'd7;
//6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd65,6'd66,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd84: Enemy_img = 4'd6;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd63,6'd64: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd75,6'd80,6'd82: Enemy_img = 4'd14;
//6'd63,6'd65,6'd70,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd64,6'd66,6'd67,6'd69,6'd70,6'd72,6'd75,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd72,6'd74: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd6;
//6'd52: Enemy_img = 4'd13;
//6'd53,6'd54,6'd55: Enemy_img = 4'd14;
//6'd56,6'd70,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53: Enemy_img = 4'd13;
//6'd51,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd57,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd6;
//6'd53: Enemy_img = 4'd13;
//6'd51,6'd56: Enemy_img = 4'd14;
//6'd35,6'd37,6'd50,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd6;
//6'd36: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd44,6'd61,6'd62,6'd63,6'd66,6'd69,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd73: Enemy_img = 4'd7;
//6'd37: Enemy_img = 4'd14;
//6'd36,6'd38,6'd39,6'd40,6'd42,6'd44,6'd45,6'd49,6'd50,6'd52,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd67,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd6;
//6'd73,6'd74: Enemy_img = 4'd7;
//6'd37,6'd38: Enemy_img = 4'd14;
//6'd39,6'd40,6'd47,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57,6'd59,6'd60,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd72,6'd73: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd36,6'd40,6'd41,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd57,6'd58,6'd60,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66,6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd73,6'd74: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39: Enemy_img = 4'd14;
//6'd36,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd52,6'd56,6'd58,6'd59,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd67,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd66,6'd72,6'd73,6'd74: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd37,6'd42,6'd43,6'd44,6'd47,6'd50,6'd55,6'd56,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd47,6'd63,6'd64,6'd76,6'd77,6'd78: Enemy_img = 4'd6;
//6'd48,6'd65,6'd66,6'd67,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd37,6'd43,6'd44,6'd50,6'd51,6'd52,6'd55,6'd56,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd63,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd6;
//6'd47,6'd48,6'd59,6'd60,6'd61,6'd62,6'd64,6'd65,6'd66,6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd70: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd46,6'd47,6'd63,6'd64,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd6;
//6'd45,6'd48,6'd59,6'd60,6'd61,6'd62,6'd65,6'd72,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd37,6'd51,6'd52,6'd55,6'd56,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd63,6'd64,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd6;
//6'd48,6'd59,6'd60,6'd61,6'd62,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd37,6'd38,6'd55,6'd56,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd45,6'd46,6'd47,6'd48,6'd63,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd44,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd38,6'd50,6'd51,6'd55,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd59,6'd60,6'd62,6'd63,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd61,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42: Enemy_img = 4'd14;
//6'd38,6'd51,6'd52,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd58,6'd59,6'd60,6'd61,6'd62,6'd64,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd49,6'd50,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd46: Enemy_img = 4'd14;
//6'd66,6'd67,6'd69,6'd70,6'd71: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd58,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd6;
//6'd54,6'd55,6'd57,6'd59,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd14;
//6'd36,6'd67,6'd68: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd50,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd35,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd68,6'd70,6'd73: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd54,6'd55,6'd57,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95: Enemy_img = 4'd6;
//6'd52,6'd53,6'd56,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd7;
//6'd34,6'd35,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd14;
//6'd38,6'd49,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd90: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd34: Enemy_img = 4'd13;
//6'd33,6'd35,6'd36,6'd46: Enemy_img = 4'd14;
//6'd37,6'd38,6'd49,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd6;
//6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87: Enemy_img = 4'd7;
//6'd35: Enemy_img = 4'd13;
//6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52: Enemy_img = 4'd6;
//6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd7;
//6'd33,6'd34,6'd35,6'd39,6'd42,6'd43,6'd46,6'd47: Enemy_img = 4'd14;
//6'd31,6'd32,6'd37,6'd38,6'd40,6'd41,6'd44,6'd45,6'd48,6'd49,6'd63,6'd91,6'd93,6'd94,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd38,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd32,6'd33,6'd37,6'd39,6'd40,6'd45,6'd46,6'd47,6'd48,6'd64,6'd65,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd60,6'd61: Enemy_img = 4'd6;
//6'd50,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd7;
//6'd35,6'd38,6'd41: Enemy_img = 4'd14;
//6'd33,6'd37,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd78,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93,6'd95,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd60,6'd61,6'd62,6'd98,6'd99: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd7;
//6'd39: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd44,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd80,6'd85,6'd87,6'd90,6'd91,6'd92,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd61,6'd98: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd50,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd7;
//6'd38,6'd41: Enemy_img = 4'd14;
//6'd36,6'd37,6'd39,6'd40,6'd42,6'd43,6'd52,6'd53,6'd65,6'd66,6'd68,6'd70,6'd72,6'd73,6'd74,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd89,6'd91,6'd92,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd57,6'd58,6'd61,6'd62,6'd98: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd56,6'd59,6'd60: Enemy_img = 4'd7;
//6'd40,6'd41: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd51,6'd53,6'd54,6'd66,6'd67,6'd69,6'd70,6'd73,6'd74,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd63: Enemy_img = 4'd7;
//6'd37,6'd38: Enemy_img = 4'd14;
//6'd36,6'd39,6'd40,6'd41,6'd42,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd67,6'd68,6'd69,6'd71,6'd72,6'd76,6'd77,6'd78,6'd79,6'd81,6'd82,6'd84,6'd85,6'd86,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd58,6'd60,6'd61,6'd62,6'd63,6'd97,6'd98: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd64: Enemy_img = 4'd7;
//6'd37,6'd38: Enemy_img = 4'd14;
//6'd36,6'd39,6'd40,6'd41,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd68,6'd69,6'd70,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd83,6'd85,6'd87,6'd88,6'd91,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd62,6'd63,6'd64,6'd65,6'd97,6'd98: Enemy_img = 4'd6;
//6'd61,6'd96: Enemy_img = 4'd7;
//6'd37,6'd38,6'd55: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd40,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd69,6'd70,6'd72,6'd73,6'd75,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd90,6'd91,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd45,6'd46,6'd49,6'd63,6'd64,6'd66,6'd97,6'd98: Enemy_img = 4'd6;
//6'd44,6'd62,6'd65: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd52,6'd56,6'd57,6'd58: Enemy_img = 4'd14;
//6'd35,6'd39,6'd50,6'd51,6'd55,6'd59,6'd69,6'd71,6'd72,6'd78,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd63,6'd97,6'd98: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd64,6'd65,6'd66,6'd67,6'd96: Enemy_img = 4'd7;
//6'd37,6'd38,6'd52,6'd56,6'd58,6'd59,6'd79: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd53,6'd55,6'd57,6'd60,6'd70,6'd71,6'd72,6'd76,6'd77,6'd78,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd64,6'd97,6'd98: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd65,6'd66,6'd67,6'd68,6'd96: Enemy_img = 4'd7;
//6'd35,6'd36,6'd37,6'd49,6'd52,6'd53,6'd59,6'd60,6'd76,6'd77,6'd78: Enemy_img = 4'd14;
//6'd34,6'd38,6'd39,6'd40,6'd46,6'd47,6'd48,6'd50,6'd51,6'd55,6'd56,6'd57,6'd58,6'd61,6'd73,6'd74,6'd75,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd97,6'd98: Enemy_img = 4'd6;
//6'd43,6'd65,6'd66,6'd95,6'd96: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd48,6'd49,6'd50,6'd51,6'd57,6'd61,6'd72,6'd74,6'd75,6'd77,6'd79: Enemy_img = 4'd14;
//6'd34,6'd35,6'd39,6'd40,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd62,6'd68,6'd71,6'd73,6'd76,6'd78,6'd80,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd66,6'd95,6'd96: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd59,6'd60,6'd61,6'd62,6'd67,6'd68,6'd70,6'd73,6'd74,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd33,6'd34,6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd56,6'd57,6'd58,6'd63,6'd69,6'd71,6'd72,6'd76,6'd77,6'd80,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd95,6'd96: Enemy_img = 4'd7;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd43,6'd46,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd60,6'd61,6'd63,6'd64,6'd68,6'd71,6'd76,6'd79: Enemy_img = 4'd14;
//6'd33,6'd34,6'd40,6'd41,6'd42,6'd44,6'd45,6'd47,6'd54,6'd55,6'd56,6'd58,6'd59,6'd62,6'd69,6'd70,6'd72,6'd75,6'd77,6'd78,6'd80,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd2;
//6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd95,6'd96: Enemy_img = 4'd7;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd58,6'd61,6'd63,6'd64,6'd65,6'd68,6'd69,6'd72,6'd75,6'd78,6'd79: Enemy_img = 4'd14;
//6'd33,6'd41,6'd45,6'd54,6'd55,6'd56,6'd59,6'd60,6'd62,6'd70,6'd71,6'd76,6'd77,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd96,6'd97: Enemy_img = 4'd7;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd57,6'd60,6'd61,6'd62,6'd64,6'd65,6'd67,6'd68,6'd69,6'd70,6'd75,6'd76,6'd79,6'd80: Enemy_img = 4'd14;
//6'd32,6'd46,6'd54,6'd56,6'd58,6'd59,6'd63,6'd71,6'd72,6'd77,6'd78,6'd84,6'd87,6'd88,6'd89,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd40,6'd42,6'd43,6'd45,6'd46,6'd96,6'd97: Enemy_img = 4'd7;
//6'd32,6'd34,6'd35,6'd36,6'd37,6'd48,6'd50,6'd51,6'd52,6'd53,6'd57,6'd60,6'd61,6'd62,6'd63,6'd65,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd80: Enemy_img = 4'd14;
//6'd31,6'd33,6'd54,6'd56,6'd58,6'd59,6'd64,6'd72,6'd78,6'd79,6'd81,6'd86,6'd88,6'd89,6'd91,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74: Enemy_img = 4'd2;
//6'd99,6'd100,6'd101: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd31,6'd34,6'd51,6'd52,6'd53,6'd57,6'd58,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd75: Enemy_img = 4'd14;
//6'd32,6'd33,6'd54,6'd55,6'd56,6'd59,6'd60,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd70,6'd73,6'd77: Enemy_img = 4'd2;
//6'd34,6'd36,6'd37,6'd38,6'd40,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd6;
//6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd30,6'd32,6'd57,6'd58,6'd59,6'd60,6'd64,6'd66,6'd67,6'd68,6'd81,6'd82: Enemy_img = 4'd14;
//6'd53,6'd55,6'd56,6'd75,6'd76,6'd79,6'd80,6'd83,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd2;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd97,6'd98,6'd99: Enemy_img = 4'd7;
//6'd63,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd56,6'd60,6'd62,6'd75,6'd76,6'd78,6'd79,6'd83,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77: Enemy_img = 4'd2;
//6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd6;
//6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd58,6'd60,6'd84,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd2;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd7;
//6'd58,6'd59,6'd60,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd55,6'd61,6'd82,6'd85,6'd86,6'd88,6'd89,6'd91,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd105,6'd106,6'd107: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd7;
//6'd57,6'd58,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd75,6'd80,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd56,6'd59,6'd60,6'd78,6'd79,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd7;
//6'd83: Enemy_img = 4'd9;
//6'd59,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd84,6'd87,6'd88: Enemy_img = 4'd14;
//6'd55,6'd56,6'd58,6'd60,6'd82,6'd85,6'd86,6'd89,6'd90,6'd93,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd7;
//6'd81,6'd82: Enemy_img = 4'd9;
//6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd85,6'd89: Enemy_img = 4'd14;
//6'd55,6'd56,6'd57,6'd61,6'd86,6'd87,6'd88,6'd95,6'd96,6'd97,6'd98,6'd110,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd80,6'd81: Enemy_img = 4'd10;
//6'd59,6'd61,6'd62,6'd64,6'd65,6'd68,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd84,6'd85,6'd86,6'd88: Enemy_img = 4'd14;
//6'd56,6'd60,6'd87,6'd89,6'd90,6'd94,6'd95,6'd96,6'd97,6'd106,6'd108,6'd109,6'd110,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd77,6'd79: Enemy_img = 4'd9;
//6'd80: Enemy_img = 4'd10;
//6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd14;
//6'd56,6'd57,6'd60,6'd83,6'd87,6'd93,6'd94,6'd95,6'd96,6'd98,6'd100,6'd101,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd78,6'd79: Enemy_img = 4'd9;
//6'd57,6'd59,6'd60,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd74,6'd75,6'd82,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd55,6'd56,6'd61,6'd63,6'd64,6'd83,6'd84,6'd88,6'd89,6'd93,6'd94,6'd95,6'd96,6'd97,6'd100,6'd101,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd57,6'd61,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd72,6'd74,6'd76,6'd78,6'd79,6'd81,6'd82,6'd83,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd55,6'd56,6'd58,6'd60,6'd62,6'd63,6'd65,6'd71,6'd84,6'd85,6'd92,6'd94,6'd95,6'd96,6'd97,6'd99,6'd100,6'd101,6'd102,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51: Enemy_img = 4'd6;
//6'd52,6'd53: Enemy_img = 4'd7;
//6'd57,6'd58,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87: Enemy_img = 4'd14;
//6'd56,6'd66,6'd70,6'd85,6'd86,6'd88,6'd89,6'd91,6'd92,6'd93,6'd95,6'd96,6'd100,6'd101,6'd102,6'd103,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52: Enemy_img = 4'd6;
//6'd53,6'd54: Enemy_img = 4'd7;
//6'd57,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd14;
//6'd55,6'd56,6'd58,6'd59,6'd67,6'd69,6'd86,6'd87,6'd88,6'd91,6'd92,6'd93,6'd94,6'd97,6'd99,6'd100,6'd101,6'd102,6'd103,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd89,6'd91: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54: Enemy_img = 4'd7;
//6'd57,6'd58,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd55,6'd56,6'd62,6'd68,6'd74,6'd87,6'd93,6'd94,6'd95,6'd97,6'd100,6'd101,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd6;
//6'd53: Enemy_img = 4'd7;
//6'd57,6'd58,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd56,6'd59,6'd61,6'd62,6'd63,6'd67,6'd73,6'd74,6'd75,6'd94,6'd95,6'd96,6'd98,6'd99,6'd102,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd87,6'd88,6'd92,6'd93: Enemy_img = 4'd6;
//6'd53,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd57,6'd58,6'd59,6'd62,6'd63,6'd65,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85: Enemy_img = 4'd14;
//6'd55,6'd56,6'd61,6'd64,6'd66,6'd67,6'd72,6'd75,6'd95,6'd96,6'd99,6'd100,6'd101,6'd102,6'd103,6'd105,6'd106,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd88,6'd93,6'd94: Enemy_img = 4'd6;
//6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd56,6'd58,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd74,6'd75,6'd78,6'd79,6'd81,6'd85: Enemy_img = 4'd14;
//6'd55,6'd57,6'd59,6'd60,6'd65,6'd68,6'd71,6'd72,6'd73,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd87,6'd88,6'd93,6'd94: Enemy_img = 4'd6;
//6'd89,6'd90,6'd91,6'd92,6'd95: Enemy_img = 4'd7;
//6'd55,6'd56,6'd57,6'd59,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd75,6'd76,6'd77,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd54,6'd58,6'd60,6'd64,6'd69,6'd70,6'd73,6'd74,6'd97,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd88,6'd89,6'd94: Enemy_img = 4'd6;
//6'd90,6'd91,6'd92,6'd93,6'd95,6'd96: Enemy_img = 4'd7;
//6'd56,6'd59,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86: Enemy_img = 4'd14;
//6'd54,6'd55,6'd57,6'd58,6'd60,6'd73,6'd98,6'd99,6'd100,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd92,6'd96,6'd97: Enemy_img = 4'd7;
//6'd55,6'd58,6'd59,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd54,6'd56,6'd57,6'd60,6'd61,6'd62,6'd63,6'd72,6'd79,6'd99,6'd100,6'd101,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd55,6'd58,6'd61,6'd62,6'd64,6'd70,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd54,6'd56,6'd57,6'd59,6'd60,6'd63,6'd65,6'd72,6'd78,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd93,6'd94,6'd95,6'd96,6'd97,6'd99: Enemy_img = 4'd6;
//6'd67,6'd68,6'd69,6'd70,6'd91,6'd92,6'd98: Enemy_img = 4'd7;
//6'd54,6'd55,6'd60,6'd61,6'd62,6'd63,6'd74,6'd76,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd53,6'd56,6'd57,6'd58,6'd59,6'd78,6'd79,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd95,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd54,6'd56,6'd57,6'd61,6'd77,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd53,6'd55,6'd58,6'd59,6'd78,6'd79,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd95,6'd96,6'd99,6'd100,6'd101: Enemy_img = 4'd6;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd93,6'd94,6'd97,6'd98: Enemy_img = 4'd7;
//6'd54,6'd56,6'd57,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91: Enemy_img = 4'd14;
//6'd52,6'd53,6'd55,6'd79,6'd80,6'd103,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd96,6'd101: Enemy_img = 4'd6;
//6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd53,6'd54,6'd80,6'd81,6'd82,6'd83,6'd84,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd61,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd75,6'd76,6'd77,6'd78,6'd79,6'd98,6'd99: Enemy_img = 4'd7;
//6'd52,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd72,6'd73,6'd74,6'd75,6'd96,6'd97: Enemy_img = 4'd6;
//6'd76,6'd77,6'd78,6'd79,6'd80,6'd98: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd74,6'd75,6'd76,6'd97,6'd98: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd14;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75,6'd76: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd81,6'd82: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd76,6'd77: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77: Enemy_img = 4'd6;
//6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97: Enemy_img = 4'd14;
//6'd96,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78: Enemy_img = 4'd6;
//6'd79: Enemy_img = 4'd7;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93: Enemy_img = 4'd14;
//6'd81,6'd92,6'd94,6'd96,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78: Enemy_img = 4'd6;
//6'd79: Enemy_img = 4'd7;
//6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd78: Enemy_img = 4'd6;
//6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd14;
//6'd80,6'd81,6'd89,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82,6'd83,6'd84,6'd85,6'd87: Enemy_img = 4'd14;
//6'd80,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd81,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd80,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80,6'd81,6'd82: Enemy_img = 4'd14;
//6'd79,6'd83,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd80: Enemy_img = 4'd14;
//6'd79,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61: Enemy_img = 4'd6;
//6'd58: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62: Enemy_img = 4'd6;
//6'd57,6'd58,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd56,6'd57,6'd59: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd42,6'd53,6'd54,6'd55,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd6;
//6'd62,6'd63: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd52,6'd54,6'd55,6'd58,6'd59,6'd60: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd66,6'd67,6'd68: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd7;
//6'd41,6'd42: Enemy_img = 4'd14;
//6'd43,6'd44,6'd52,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69,6'd70: Enemy_img = 4'd6;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd14;
//6'd45,6'd50,6'd51,6'd52,6'd59,6'd60,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd83,6'd85,6'd87: Enemy_img = 4'd6;
//6'd63,6'd64,6'd65: Enemy_img = 4'd7;
//6'd40,6'd41: Enemy_img = 4'd13;
//6'd42,6'd43: Enemy_img = 4'd14;
//6'd49,6'd50,6'd51,6'd59,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd7;
//6'd42: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41: Enemy_img = 4'd14;
//6'd49,6'd61,6'd88,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84: Enemy_img = 4'd6;
//6'd56,6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd7;
//6'd39,6'd40: Enemy_img = 4'd14;
//6'd46,6'd47,6'd50,6'd61,6'd62,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd92: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd80,6'd81,6'd82: Enemy_img = 4'd7;
//6'd39,6'd44,6'd45,6'd47,6'd48,6'd60,6'd61,6'd86,6'd87,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd75,6'd92: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd45,6'd49,6'd61,6'd62,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd92: Enemy_img = 4'd6;
//6'd53,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd43,6'd46,6'd47,6'd62,6'd63,6'd64,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd93: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78: Enemy_img = 4'd7;
//6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd46,6'd47,6'd61,6'd62,6'd63,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd92,6'd93: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75: Enemy_img = 4'd7;
//6'd27,6'd29,6'd30,6'd31,6'd33,6'd35,6'd37,6'd38,6'd39,6'd46,6'd47,6'd48,6'd59,6'd62,6'd64,6'd66,6'd81,6'd82,6'd85,6'd86,6'd87,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd93,6'd94: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd37,6'd38,6'd39,6'd41,6'd42,6'd44,6'd46,6'd47,6'd59,6'd60,6'd66,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd88,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57,6'd93,6'd94: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd69,6'd70,6'd92: Enemy_img = 4'd7;
//6'd27,6'd28,6'd29: Enemy_img = 4'd14;
//6'd26,6'd30,6'd31,6'd34,6'd38,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd61,6'd63,6'd64,6'd65,6'd66,6'd67,6'd77,6'd80,6'd82,6'd89,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd52,6'd53,6'd54,6'd93,6'd94: Enemy_img = 4'd6;
//6'd40,6'd92: Enemy_img = 4'd7;
//6'd28,6'd29,6'd30,6'd31: Enemy_img = 4'd14;
//6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd44,6'd48,6'd63,6'd64,6'd65,6'd66,6'd90,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd52,6'd53,6'd94,6'd95: Enemy_img = 4'd6;
//6'd40,6'd41,6'd93: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd33,6'd34: Enemy_img = 4'd14;
//6'd28,6'd32,6'd35,6'd36,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd73,6'd75,6'd76,6'd78,6'd80,6'd81,6'd82,6'd87,6'd91: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd51,6'd52,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd38,6'd40,6'd41,6'd92,6'd93: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd28,6'd44,6'd46,6'd58,6'd70,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40,6'd41,6'd52,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd38,6'd51,6'd93: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd29,6'd45,6'd68,6'd69,6'd70,6'd72,6'd73,6'd76,6'd77,6'd78,6'd81,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd50,6'd51,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd44,6'd48,6'd93,6'd94: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd34,6'd35: Enemy_img = 4'd14;
//6'd30,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd73,6'd74,6'd75,6'd80,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48,6'd49,6'd50,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd38,6'd39,6'd40,6'd47,6'd51,6'd52,6'd93,6'd94: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Enemy_img = 4'd14;
//6'd30,6'd59,6'd61,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd46,6'd96,6'd97,6'd98: Enemy_img = 4'd6;
//6'd38,6'd39,6'd45,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd94,6'd95: Enemy_img = 4'd7;
//6'd31,6'd33,6'd34,6'd35,6'd36,6'd41: Enemy_img = 4'd14;
//6'd32,6'd60,6'd62,6'd63,6'd64,6'd65,6'd67,6'd70,6'd73,6'd74,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd94,6'd95,6'd96: Enemy_img = 4'd7;
//6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd14;
//6'd31,6'd32,6'd60,6'd66,6'd69,6'd73,6'd77,6'd80,6'd81,6'd82,6'd83,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd57,6'd58,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd6;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd95,6'd96,6'd97: Enemy_img = 4'd7;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd77: Enemy_img = 4'd14;
//6'd32,6'd44,6'd62,6'd63,6'd64,6'd66,6'd70,6'd73,6'd76,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd57,6'd58,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd107,6'd108: Enemy_img = 4'd6;
//6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd96,6'd97: Enemy_img = 4'd7;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd76: Enemy_img = 4'd14;
//6'd45,6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd74,6'd75,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd93,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd59,6'd60,6'd101,6'd102,6'd103,6'd104,6'd106,6'd109: Enemy_img = 4'd6;
//6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61,6'd97,6'd98,6'd99,6'd100,6'd105,6'd107: Enemy_img = 4'd7;
//6'd34,6'd36,6'd37,6'd38,6'd39,6'd75,6'd76,6'd78: Enemy_img = 4'd14;
//6'd32,6'd33,6'd35,6'd42,6'd44,6'd45,6'd67,6'd69,6'd70,6'd71,6'd74,6'd77,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd91,6'd92,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd58,6'd59,6'd60,6'd63: Enemy_img = 4'd6;
//6'd47,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61,6'd62,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd42,6'd43,6'd73,6'd74,6'd78,6'd79: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd40,6'd41,6'd44,6'd45,6'd67,6'd69,6'd70,6'd72,6'd75,6'd76,6'd77,6'd82,6'd83,6'd84,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd6;
//6'd53,6'd54,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd7;
//6'd31,6'd32,6'd39,6'd43,6'd73,6'd74,6'd76,6'd78,6'd79: Enemy_img = 4'd14;
//6'd37,6'd38,6'd40,6'd41,6'd42,6'd44,6'd45,6'd50,6'd69,6'd71,6'd72,6'd75,6'd77,6'd80,6'd81,6'd86,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd110,6'd111,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd56,6'd58,6'd59,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd60,6'd64,6'd65,6'd66,6'd67,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd37,6'd39,6'd40,6'd41,6'd72,6'd73,6'd74,6'd76,6'd78,6'd79,6'd80: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd38,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd70,6'd71,6'd75,6'd77,6'd81,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95,6'd96,6'd97,6'd98,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47,6'd61,6'd62,6'd63: Enemy_img = 4'd6;
//6'd64,6'd65,6'd66,6'd103: Enemy_img = 4'd7;
//6'd30,6'd31: Enemy_img = 4'd13;
//6'd32,6'd35,6'd36,6'd37,6'd39,6'd40,6'd70,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd34,6'd38,6'd41,6'd42,6'd43,6'd49,6'd52,6'd53,6'd54,6'd55,6'd57,6'd68,6'd69,6'd71,6'd72,6'd77,6'd78,6'd82,6'd83,6'd87,6'd88,6'd90,6'd95,6'd96,6'd97,6'd99,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74: Enemy_img = 4'd2;
//6'd47,6'd63,6'd64: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd65: Enemy_img = 4'd7;
//6'd32,6'd33: Enemy_img = 4'd13;
//6'd30,6'd31,6'd36,6'd38,6'd39,6'd54,6'd57,6'd67,6'd68,6'd71,6'd72,6'd73,6'd76,6'd77,6'd83: Enemy_img = 4'd14;
//6'd35,6'd37,6'd40,6'd42,6'd49,6'd50,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60,6'd69,6'd70,6'd79,6'd80,6'd81,6'd82,6'd84,6'd91,6'd92,6'd95,6'd96,6'd99,6'd100,6'd104,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75: Enemy_img = 4'd2;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd66: Enemy_img = 4'd7;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd55,6'd56,6'd58,6'd59,6'd68,6'd69,6'd70,6'd76,6'd77,6'd80,6'd82,6'd83,6'd91,6'd92: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd50,6'd51,6'd52,6'd53,6'd54,6'd57,6'd60,6'd61,6'd62,6'd71,6'd72,6'd73,6'd81,6'd84,6'd85,6'd86,6'd90,6'd93,6'd95,6'd97,6'd98,6'd99,6'd100,6'd103,6'd104,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd79: Enemy_img = 4'd2;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd32,6'd33,6'd37,6'd40,6'd51,6'd56,6'd61,6'd62,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72,6'd76,6'd82,6'd83,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd29,6'd30,6'd31,6'd35,6'd36,6'd38,6'd39,6'd41,6'd50,6'd52,6'd55,6'd57,6'd58,6'd59,6'd60,6'd63,6'd73,6'd77,6'd81,6'd86,6'd87,6'd91,6'd92,6'd93,6'd97,6'd98,6'd99,6'd103,6'd104,6'd105,6'd106,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd75,6'd79: Enemy_img = 4'd2;
//6'd48,6'd49: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd37,6'd39,6'd40,6'd58,6'd61,6'd62,6'd64,6'd65,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd81,6'd82,6'd83,6'd89,6'd90,6'd92: Enemy_img = 4'd14;
//6'd31,6'd32,6'd35,6'd36,6'd38,6'd41,6'd50,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd59,6'd60,6'd63,6'd77,6'd85,6'd87,6'd88,6'd91,6'd93,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd103,6'd104,6'd105,6'd106,6'd107,6'd109,6'd110,6'd111,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd73,6'd80: Enemy_img = 4'd2;
//6'd45,6'd46,6'd47,6'd49: Enemy_img = 4'd6;
//6'd44: Enemy_img = 4'd7;
//6'd39,6'd52,6'd53,6'd57,6'd60,6'd61,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd77,6'd81,6'd82,6'd83,6'd87,6'd88,6'd92: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd51,6'd54,6'd56,6'd58,6'd59,6'd63,6'd64,6'd78,6'd85,6'd89,6'd90,6'd91,6'd93,6'd96,6'd97,6'd98,6'd99,6'd100,6'd104,6'd105,6'd106,6'd107,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd79,6'd80: Enemy_img = 4'd2;
//6'd43,6'd44,6'd45: Enemy_img = 4'd6;
//6'd85,6'd86: Enemy_img = 4'd9;
//6'd37,6'd38,6'd51,6'd58,6'd59,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd74,6'd75,6'd76,6'd83,6'd88,6'd89,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd39,6'd41,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd57,6'd60,6'd61,6'd65,6'd82,6'd90,6'd93,6'd99,6'd100,6'd104,6'd105,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd77,6'd78: Enemy_img = 4'd2;
//6'd41,6'd42: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45: Enemy_img = 4'd7;
//6'd84,6'd86: Enemy_img = 4'd9;
//6'd85: Enemy_img = 4'd10;
//6'd37,6'd38,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd81,6'd82,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd36,6'd39,6'd40,6'd47,6'd48,6'd49,6'd55,6'd57,6'd61,6'd91,6'd92,6'd93,6'd96,6'd97,6'd98,6'd102,6'd107,6'd108,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43: Enemy_img = 4'd6;
//6'd44,6'd45: Enemy_img = 4'd7;
//6'd84,6'd85: Enemy_img = 4'd10;
//6'd37,6'd38,6'd39,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd62,6'd63,6'd64,6'd65,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd79,6'd80,6'd81,6'd82,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd40,6'd47,6'd48,6'd56,6'd57,6'd58,6'd60,6'd61,6'd87,6'd93,6'd96,6'd97,6'd98,6'd99,6'd100,6'd104,6'd105,6'd107,6'd108,6'd109,6'd110,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd42,6'd43: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd84: Enemy_img = 4'd9;
//6'd85: Enemy_img = 4'd10;
//6'd37,6'd38,6'd39,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd63,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd87,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd40,6'd48,6'd56,6'd58,6'd62,6'd65,6'd88,6'd89,6'd93,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd96,6'd97: Enemy_img = 4'd6;
//6'd83,6'd84: Enemy_img = 4'd9;
//6'd38,6'd39,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd59,6'd60,6'd61,6'd62,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd36,6'd37,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd56,6'd58,6'd65,6'd90,6'd91,6'd92,6'd93,6'd101,6'd102,6'd104,6'd105,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd82,6'd83: Enemy_img = 4'd9;
//6'd37,6'd38,6'd39,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd60,6'd61,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd57,6'd59,6'd63,6'd93,6'd103,6'd104,6'd105,6'd106,6'd107,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd100,6'd101: Enemy_img = 4'd6;
//6'd95,6'd96,6'd97,6'd98,6'd99,6'd102: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd46,6'd47,6'd51,6'd53,6'd54,6'd63,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd48,6'd49,6'd56,6'd59,6'd60,6'd62,6'd64,6'd65,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd100,6'd101,6'd102: Enemy_img = 4'd6;
//6'd49,6'd52,6'd55,6'd57,6'd95,6'd96,6'd97,6'd98,6'd99,6'd103,6'd104: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd62,6'd63,6'd64,6'd66,6'd67,6'd69,6'd70,6'd71,6'd73,6'd75,6'd76,6'd79,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd36,6'd37,6'd44,6'd61,6'd65,6'd108,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd95,6'd96,6'd101,6'd102,6'd107: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd97,6'd98,6'd99,6'd100,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd62,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd60,6'd63,6'd64,6'd65,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95,6'd96,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd97,6'd100: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd64,6'd65,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93: Enemy_img = 4'd14;
//6'd36,6'd37,6'd60,6'd61,6'd63,6'd66,6'd77,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd110: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd109: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd14;
//6'd36,6'd60,6'd61,6'd62,6'd66,6'd70,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd51,6'd99,6'd104,6'd105: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd100,6'd101,6'd102,6'd103,6'd106,6'd107,6'd108: Enemy_img = 4'd7;
//6'd37,6'd38,6'd39,6'd40,6'd68,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd14;
//6'd36,6'd61,6'd62,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd76,6'd80,6'd81,6'd82,6'd83: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd104,6'd105,6'd106: Enemy_img = 4'd6;
//6'd42,6'd55,6'd56,6'd57,6'd58,6'd59,6'd102,6'd103,6'd107,6'd108: Enemy_img = 4'd7;
//6'd39,6'd65,6'd66,6'd70,6'd71,6'd72,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd85,6'd86,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd61,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd105,6'd106,6'd107: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd104,6'd108: Enemy_img = 4'd7;
//6'd36,6'd63,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101: Enemy_img = 4'd14;
//6'd37,6'd62,6'd64,6'd66,6'd67,6'd75,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd41,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd107,6'd108: Enemy_img = 4'd6;
//6'd57,6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd7;
//6'd36,6'd37,6'd64,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd78,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd62,6'd63,6'd65,6'd75,6'd79,6'd80,6'd81,6'd82,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61: Enemy_img = 4'd7;
//6'd35,6'd65,6'd68,6'd69,6'd72,6'd73,6'd78,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd62,6'd63,6'd64,6'd66,6'd70,6'd71,6'd74,6'd75,6'd76,6'd77,6'd79,6'd82,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61: Enemy_img = 4'd7;
//6'd64,6'd65,6'd66,6'd71,6'd75,6'd76,6'd79,6'd80,6'd83,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd63,6'd70,6'd72,6'd73,6'd74,6'd77,6'd78,6'd81,6'd82,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd65,6'd66,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd90,6'd91,6'd92,6'd93,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//6'd64,6'd67,6'd68,6'd69,6'd73,6'd74,6'd88,6'd89,6'd108,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd61,6'd62: Enemy_img = 4'd7;
//6'd65,6'd66,6'd67,6'd68,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd87,6'd90,6'd91,6'd92,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//6'd64,6'd73,6'd82,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd61,6'd62,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd7;
//6'd66,6'd67,6'd68,6'd72,6'd74,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd64,6'd65,6'd69,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd69,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd64,6'd65,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd93,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62,6'd80,6'd81,6'd83,6'd85,6'd86: Enemy_img = 4'd6;
//6'd77,6'd78,6'd79,6'd82,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd7;
//6'd65,6'd66,6'd69,6'd70,6'd72,6'd73,6'd74,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd64,6'd67,6'd68,6'd71,6'd93,6'd94,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd76,6'd77,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd7;
//6'd66,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd14;
//6'd64,6'd65,6'd67,6'd70,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd74,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd66,6'd68,6'd69,6'd71,6'd72,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd64,6'd65,6'd67,6'd70,6'd94,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd74,6'd75,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd6;
//6'd91,6'd92: Enemy_img = 4'd7;
//6'd65,6'd66,6'd71,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd14;
//6'd67,6'd68,6'd69,6'd70,6'd94,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd72,6'd73,6'd74,6'd75,6'd76,6'd89,6'd90: Enemy_img = 4'd6;
//6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd66,6'd68,6'd69,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd65,6'd67,6'd70,6'd94,6'd100,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd71,6'd72,6'd73,6'd91: Enemy_img = 4'd6;
//6'd92,6'd93: Enemy_img = 4'd7;
//6'd65,6'd68,6'd69,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd66,6'd67,6'd95,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd91,6'd92: Enemy_img = 4'd6;
//6'd66,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd14;
//6'd65,6'd67,6'd94,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd93: Enemy_img = 4'd6;
//6'd66,6'd67,6'd96,6'd97: Enemy_img = 4'd14;
//6'd65,6'd95,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65,6'd96: Enemy_img = 4'd14;
//6'd94,6'd95,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd65: Enemy_img = 4'd14;
//6'd95,6'd96: Enemy_img = 4'd15;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd6;
//6'd43,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd79: Enemy_img = 4'd6;
//6'd43,6'd44,6'd75,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd70,6'd71,6'd72,6'd80: Enemy_img = 4'd6;
//6'd43,6'd77,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd68,6'd69,6'd70,6'd71,6'd80,6'd81: Enemy_img = 4'd6;
//6'd43,6'd45,6'd74,6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd66,6'd67,6'd68,6'd69,6'd70,6'd81,6'd82: Enemy_img = 4'd6;
//6'd45,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd48,6'd69,6'd70: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd48,6'd49,6'd68,6'd69: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd73,6'd74,6'd75,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd66,6'd67,6'd68,6'd69,6'd82: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd65,6'd66,6'd67,6'd68,6'd83: Enemy_img = 4'd7;
//6'd44,6'd46,6'd47,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd83,6'd84: Enemy_img = 4'd7;
//6'd41,6'd42,6'd46,6'd47,6'd48,6'd71,6'd72,6'd74,6'd81,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88,6'd89,6'd90,6'd99,6'd100,6'd101: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd84,6'd85: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd47,6'd48,6'd70,6'd71,6'd72,6'd77,6'd78,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd84,6'd85,6'd86,6'd100: Enemy_img = 4'd7;
//6'd40,6'd42,6'd43,6'd48,6'd50,6'd69,6'd70,6'd78,6'd79,6'd80,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd85,6'd86,6'd87,6'd88,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd40,6'd50,6'd51,6'd68,6'd73,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd86,6'd87,6'd88,6'd89,6'd90,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd50,6'd51,6'd52,6'd71,6'd72,6'd73,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd6;
//6'd46,6'd47,6'd58,6'd59,6'd60,6'd61,6'd62,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd39,6'd40,6'd51,6'd52,6'd53,6'd54,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd60,6'd61,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd52,6'd53,6'd54,6'd55,6'd57,6'd67,6'd68,6'd69,6'd70,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd86,6'd87,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd6;
//6'd46,6'd47,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34: Enemy_img = 4'd14;
//6'd39,6'd40,6'd52,6'd53,6'd57,6'd58,6'd65,6'd67,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd83,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd14;
//6'd37,6'd50,6'd55,6'd56,6'd57,6'd58,6'd65,6'd72,6'd73,6'd74,6'd75,6'd76,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd99,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd6;
//6'd44,6'd45: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32: Enemy_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd51,6'd52,6'd53,6'd55,6'd56,6'd57,6'd62,6'd65,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd94,6'd95,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd30,6'd31: Enemy_img = 4'd14;
//6'd35,6'd36,6'd55,6'd56,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd71,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87,6'd89,6'd90,6'd91,6'd94,6'd95,6'd97,6'd99,6'd100,6'd101,6'd102,6'd103,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd30,6'd31: Enemy_img = 4'd14;
//6'd36,6'd38,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd71,6'd72,6'd75,6'd76,6'd77,6'd78,6'd79,6'd85,6'd86,6'd90,6'd91,6'd93,6'd94,6'd95,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd71: Enemy_img = 4'd14;
//6'd30,6'd33,6'd38,6'd39,6'd52,6'd53,6'd59,6'd61,6'd62,6'd63,6'd64,6'd67,6'd70,6'd72,6'd73,6'd77,6'd78,6'd79,6'd81,6'd82,6'd83,6'd84,6'd85,6'd88,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd100,6'd101,6'd102,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd6;
//6'd44,6'd45: Enemy_img = 4'd7;
//6'd71,6'd73,6'd88: Enemy_img = 4'd14;
//6'd32,6'd33,6'd35,6'd38,6'd39,6'd40,6'd51,6'd58,6'd59,6'd67,6'd70,6'd72,6'd74,6'd81,6'd82,6'd83,6'd84,6'd87,6'd89,6'd93,6'd94,6'd95,6'd96,6'd97,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd70,6'd71,6'd73,6'd74,6'd87: Enemy_img = 4'd14;
//6'd31,6'd32,6'd33,6'd35,6'd39,6'd40,6'd41,6'd57,6'd58,6'd59,6'd61,6'd63,6'd64,6'd65,6'd69,6'd72,6'd75,6'd76,6'd86,6'd88,6'd89,6'd93,6'd94,6'd95,6'd96,6'd97,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45: Enemy_img = 4'd6;
//6'd46: Enemy_img = 4'd7;
//6'd74,6'd75,6'd76,6'd86,6'd87,6'd89: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd37,6'd40,6'd41,6'd55,6'd56,6'd57,6'd58,6'd59,6'd61,6'd65,6'd69,6'd70,6'd71,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd85,6'd88,6'd90,6'd109,6'd110,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd69,6'd70,6'd72,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd85,6'd86,6'd87,6'd89: Enemy_img = 4'd14;
//6'd28,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd71,6'd73,6'd78,6'd81,6'd82,6'd83,6'd84,6'd88,6'd90,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd6;
//6'd45: Enemy_img = 4'd7;
//6'd69,6'd70,6'd72,6'd79,6'd80,6'd89,6'd90: Enemy_img = 4'd14;
//6'd27,6'd28,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd38,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd65,6'd66,6'd68,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd84,6'd85,6'd86,6'd87,6'd88,6'd91,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd34,6'd44,6'd47: Enemy_img = 4'd7;
//6'd68,6'd69,6'd72,6'd73,6'd74,6'd77,6'd79,6'd80,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd26,6'd30,6'd31,6'd32,6'd36,6'd40,6'd63,6'd65,6'd67,6'd78,6'd82,6'd83,6'd88,6'd89,6'd90,6'd91,6'd94: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd76: Enemy_img = 4'd2;
//6'd33,6'd44,6'd45,6'd52,6'd53,6'd54,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd6;
//6'd34,6'd35,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd7;
//6'd84: Enemy_img = 4'd9;
//6'd73,6'd74,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd24,6'd26,6'd28,6'd38,6'd39,6'd40,6'd67,6'd68,6'd69,6'd78,6'd83,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd77: Enemy_img = 4'd2;
//6'd32,6'd33,6'd34,6'd43,6'd44,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd94,6'd95,6'd96,6'd99,6'd100,6'd101,6'd102,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd6;
//6'd35,6'd36,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd63,6'd64,6'd97,6'd98,6'd103,6'd104,6'd109: Enemy_img = 4'd7;
//6'd83,6'd84: Enemy_img = 4'd9;
//6'd67,6'd68,6'd69,6'd70,6'd74,6'd79,6'd80,6'd81,6'd87,6'd88,6'd89,6'd90,6'd91: Enemy_img = 4'd14;
//6'd23,6'd24,6'd28,6'd29,6'd30,6'd66,6'd75,6'd86,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd78: Enemy_img = 4'd2;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd94,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd6;
//6'd33,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd61,6'd62,6'd63,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd107,6'd108,6'd109: Enemy_img = 4'd7;
//6'd83: Enemy_img = 4'd9;
//6'd84: Enemy_img = 4'd10;
//6'd81: Enemy_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd80,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73,6'd78: Enemy_img = 4'd2;
//6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd42,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd94,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd6;
//6'd33,6'd37,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd61,6'd62,6'd63,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd107,6'd108,6'd109: Enemy_img = 4'd7;
//6'd83,6'd84: Enemy_img = 4'd10;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd75,6'd76,6'd80,6'd81,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd19,6'd20,6'd27: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd77: Enemy_img = 4'd2;
//6'd32,6'd33,6'd34,6'd43,6'd44,6'd53,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd62,6'd94,6'd95,6'd96,6'd99,6'd100,6'd101,6'd102,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd6;
//6'd35,6'd36,6'd42,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57,6'd58,6'd63,6'd64,6'd97,6'd98,6'd103,6'd104,6'd109: Enemy_img = 4'd7;
//6'd83: Enemy_img = 4'd9;
//6'd84: Enemy_img = 4'd10;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd66,6'd67,6'd68,6'd69,6'd70,6'd74,6'd75,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd21,6'd22: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71,6'd76: Enemy_img = 4'd2;
//6'd33,6'd44,6'd45,6'd52,6'd53,6'd54,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd6;
//6'd34,6'd35,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd7;
//6'd83,6'd84: Enemy_img = 4'd9;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38,6'd39,6'd40,6'd67,6'd68,6'd69,6'd73,6'd74,6'd78,6'd79,6'd80,6'd81,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92: Enemy_img = 4'd14;
//6'd23,6'd41: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd34,6'd44,6'd47: Enemy_img = 4'd7;
//6'd82,6'd83: Enemy_img = 4'd9;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd36,6'd37,6'd38,6'd39,6'd40,6'd63,6'd64,6'd65,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94: Enemy_img = 4'd14;
//6'd24,6'd25,6'd42,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd34,6'd40,6'd44,6'd47,6'd67,6'd81,6'd82,6'd83,6'd92,6'd101,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd46: Enemy_img = 4'd6;
//6'd45: Enemy_img = 4'd7;
//default: Enemy_img = 4'd14;
//6'd26,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd62,6'd112,6'd113: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd39,6'd44,6'd47,6'd48,6'd49,6'd67,6'd91,6'd101,6'd113,6'd114,6'd115,6'd116,6'd117,6'd118,6'd119,6'd120,6'd121,6'd122,6'd123,6'd124,6'd125,6'd126,6'd127,6'd128: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//default: Enemy_img = 4'd14;
//6'd27,6'd29,6'd40,6'd42,6'd43,6'd50,6'd51,6'd52,6'd56,6'd57,6'd58,6'd59,6'd62,6'd63,6'd64,6'd65,6'd111,6'd112: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45: Enemy_img = 4'd6;
//6'd46: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd55,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110: Enemy_img = 4'd14;
//6'd28,6'd29,6'd39,6'd42,6'd43,6'd48,6'd49,6'd52,6'd53,6'd54,6'd56,6'd58,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd57,6'd62,6'd63,6'd64,6'd65,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd30,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd51,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd6;
//6'd44,6'd45: Enemy_img = 4'd7;
//6'd32,6'd34,6'd35,6'd38,6'd39,6'd40,6'd51,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd31,6'd33,6'd37,6'd41,6'd42,6'd49,6'd50,6'd52,6'd53,6'd56,6'd57,6'd61,6'd66,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd38,6'd39,6'd52,6'd53,6'd59,6'd60,6'd64,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd86,6'd88,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd30,6'd32,6'd33,6'd36,6'd37,6'd40,6'd41,6'd50,6'd51,6'd54,6'd55,6'd57,6'd58,6'd61,6'd62,6'd63,6'd66,6'd79,6'd83,6'd84,6'd85,6'd91,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49: Enemy_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Enemy_img = 4'd7;
//6'd36,6'd38,6'd55,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd69,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd30,6'd31,6'd34,6'd35,6'd37,6'd39,6'd40,6'd51,6'd52,6'd53,6'd54,6'd56,6'd58,6'd59,6'd65,6'd79,6'd83,6'd91,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Enemy_img = 4'd7;
//6'd30,6'd31,6'd35,6'd36,6'd38,6'd39,6'd52,6'd53,6'd54,6'd55,6'd56,6'd61,6'd62,6'd63,6'd68,6'd69,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd93,6'd94,6'd95,6'd96,6'd97,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd33,6'd34,6'd37,6'd40,6'd41,6'd50,6'd51,6'd57,6'd59,6'd60,6'd65,6'd66,6'd67,6'd79,6'd83,6'd91,6'd92,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd47: Enemy_img = 4'd6;
//6'd44,6'd45: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd36,6'd40,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd62,6'd65,6'd66,6'd68,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd87,6'd88,6'd89,6'd90,6'd91,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//6'd34,6'd35,6'd37,6'd38,6'd39,6'd41,6'd42,6'd49,6'd50,6'd58,6'd60,6'd61,6'd64,6'd67,6'd79,6'd83,6'd84,6'd85,6'd86,6'd92,6'd93,6'd94,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd30,6'd31,6'd32,6'd33: Enemy_img = 4'd13;
//6'd37,6'd38,6'd40,6'd41,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd65,6'd70,6'd71,6'd72,6'd80,6'd81,6'd82,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd42,6'd43,6'd48,6'd49,6'd59,6'd61,6'd62,6'd64,6'd66,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd83,6'd86,6'd98,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd6;
//6'd46,6'd47,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd40,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd84,6'd85,6'd87,6'd88,6'd89,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: Enemy_img = 4'd14;
//6'd36,6'd37,6'd39,6'd41,6'd42,6'd49,6'd50,6'd59,6'd66,6'd69,6'd73,6'd79,6'd83,6'd86,6'd99,6'd108: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44: Enemy_img = 4'd6;
//6'd45,6'd46,6'd47,6'd48,6'd60,6'd61,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98: Enemy_img = 4'd7;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd67,6'd68,6'd74,6'd75,6'd76,6'd77,6'd78,6'd84,6'd85,6'd86,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd50,6'd51,6'd63,6'd64,6'd69,6'd70,6'd71,6'd72,6'd73,6'd79,6'd80,6'd81,6'd82,6'd83,6'd87,6'd100,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45: Enemy_img = 4'd6;
//6'd46,6'd47,6'd58,6'd59,6'd60,6'd61,6'd62,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd7;
//6'd39,6'd40,6'd51,6'd52,6'd53,6'd54,6'd69,6'd70,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd37,6'd38,6'd41,6'd42,6'd49,6'd50,6'd64,6'd65,6'd66,6'd71,6'd79,6'd101,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd86,6'd87,6'd88,6'd89,6'd90,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd72,6'd73,6'd74,6'd80,6'd81,6'd82,6'd83,6'd84,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd14;
//6'd38,6'd42,6'd43,6'd48,6'd49,6'd50,6'd51,6'd52,6'd65,6'd66,6'd67,6'd68,6'd71,6'd75,6'd76,6'd77,6'd78,6'd79,6'd101,6'd107: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd85,6'd86,6'd87,6'd88,6'd98,6'd99,6'd100: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd49,6'd50,6'd51,6'd68,6'd73,6'd74,6'd76,6'd77,6'd78,6'd80,6'd81,6'd82,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd38,6'd39,6'd43,6'd44,6'd47,6'd48,6'd66,6'd67,6'd69,6'd70,6'd75,6'd79,6'd102,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd84,6'd85,6'd86,6'd100: Enemy_img = 4'd7;
//6'd40,6'd41,6'd42,6'd49,6'd50,6'd69,6'd70,6'd76,6'd77,6'd78,6'd80,6'd103,6'd104,6'd105: Enemy_img = 4'd14;
//6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd67,6'd68,6'd71,6'd72,6'd75,6'd79,6'd102,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd86,6'd87,6'd88,6'd89,6'd90,6'd99,6'd100,6'd101: Enemy_img = 4'd6;
//6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd84,6'd85: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd47,6'd49,6'd70,6'd71,6'd72,6'd77,6'd78,6'd104: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd45,6'd46,6'd48,6'd68,6'd69,6'd73,6'd74,6'd81,6'd82,6'd103,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56,6'd57,6'd58,6'd59,6'd60,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd6;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd83,6'd84: Enemy_img = 4'd7;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd71,6'd72,6'd73,6'd74,6'd81,6'd104: Enemy_img = 4'd14;
//6'd40,6'd69,6'd70,6'd75,6'd76,6'd79,6'd80,6'd103,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd84,6'd85,6'd86: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd65,6'd66,6'd67,6'd68,6'd83: Enemy_img = 4'd7;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd81: Enemy_img = 4'd14;
//6'd40,6'd41,6'd70,6'd71,6'd77,6'd78,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd49,6'd50,6'd51,6'd66,6'd67,6'd68,6'd69,6'd82: Enemy_img = 4'd7;
//6'd44,6'd45,6'd46,6'd47,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd71,6'd72,6'd73,6'd74,6'd75,6'd78,6'd104: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd82,6'd83,6'd84: Enemy_img = 4'd6;
//6'd48,6'd49,6'd68,6'd69: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd73,6'd74,6'd76,6'd77,6'd79,6'd80: Enemy_img = 4'd14;
//6'd41,6'd42,6'd71,6'd72,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd81,6'd82,6'd83: Enemy_img = 4'd6;
//6'd48,6'd69,6'd70: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd46,6'd73,6'd74,6'd76,6'd77,6'd79: Enemy_img = 4'd14;
//6'd41,6'd42,6'd72,6'd75,6'd78: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd66,6'd67,6'd68,6'd69,6'd70,6'd81,6'd82: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd74: Enemy_img = 4'd14;
//6'd42,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd79: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd47,6'd48,6'd68,6'd69,6'd70,6'd71,6'd80,6'd81: Enemy_img = 4'd6;
//6'd45,6'd74,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd42,6'd43,6'd44,6'd73,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd70,6'd71,6'd72,6'd80: Enemy_img = 4'd6;
//6'd43,6'd75,6'd77,6'd78: Enemy_img = 4'd14;
//6'd42,6'd44,6'd74,6'd76: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd79: Enemy_img = 4'd6;
//6'd43,6'd44,6'd75: Enemy_img = 4'd14;
//6'd74,6'd76,6'd77: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd73: Enemy_img = 4'd6;
//6'd43,6'd76,6'd77: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd76,6'd77: Enemy_img = 4'd14;
//6'd75: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76: Enemy_img = 4'd14;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//// Enemy_type_4 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd19: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd90: Enemy_img = 4'd6;
//6'd63,6'd64,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd66,6'd67,6'd88,6'd89: Enemy_img = 4'd6;
//6'd63,6'd64,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd68,6'd69,6'd70,6'd88: Enemy_img = 4'd6;
//6'd89,6'd90: Enemy_img = 4'd7;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd93,6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd69,6'd70,6'd71,6'd72,6'd73,6'd86,6'd87: Enemy_img = 4'd6;
//6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd67,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd71,6'd72,6'd73,6'd74,6'd75,6'd83,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd6;
//6'd88,6'd89: Enemy_img = 4'd7;
//6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd71,6'd86,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd7;
//6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd6;
//6'd73,6'd74,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd7;
//6'd63,6'd64,6'd68,6'd69,6'd70,6'd71,6'd92,6'd93,6'd97,6'd98,6'd99,6'd100,6'd101: Enemy_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd57,6'd58,6'd59,6'd77,6'd78,6'd80,6'd82,6'd83: Enemy_img = 4'd6;
//6'd74,6'd75,6'd76,6'd79,6'd81,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd94,6'd95,6'd97,6'd98,6'd99: Enemy_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88: Enemy_img = 4'd7;
//6'd63,6'd64,6'd65,6'd66,6'd91,6'd92,6'd93,6'd94,6'd95,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55,6'd56,6'd57: Enemy_img = 4'd6;
//6'd58,6'd59,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86: Enemy_img = 4'd7;
//6'd62,6'd64,6'd65,6'd69,6'd71,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd6;
//6'd58,6'd59: Enemy_img = 4'd7;
//6'd65,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd75,6'd76,6'd77,6'd79,6'd84,6'd87,6'd90,6'd92,6'd93,6'd94,6'd95,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd55: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58,6'd59: Enemy_img = 4'd7;
//6'd62,6'd63,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd85,6'd87,6'd88,6'd93,6'd94,6'd98,6'd99,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58: Enemy_img = 4'd7;
//6'd61,6'd62,6'd63,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd80,6'd81,6'd82,6'd83,6'd84,6'd87,6'd88,6'd90,6'd95,6'd96,6'd97,6'd101,6'd102,6'd103,6'd104,6'd105: Enemy_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Enemy_img = 4'd6;
//6'd56,6'd57,6'd58: Enemy_img = 4'd7;
//6'd32,6'd62,6'd65,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd38,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd104,6'd105: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56,6'd57,6'd58: Enemy_img = 4'd7;
//6'd33,6'd34,6'd61,6'd64,6'd65,6'd67,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd78,6'd79,6'd80,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90,6'd91,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd102,6'd103,6'd104: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd57,6'd101,6'd105: Enemy_img = 4'd7;
//6'd33,6'd60,6'd63,6'd64,6'd65,6'd66,6'd68,6'd69,6'd71,6'd75,6'd76,6'd77,6'd79,6'd80,6'd87,6'd88,6'd89,6'd90,6'd93,6'd94,6'd95,6'd97,6'd98: Enemy_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd101,6'd102,6'd103: Enemy_img = 4'd6;
//6'd39,6'd52,6'd53,6'd54,6'd55,6'd56,6'd99,6'd100,6'd104,6'd105: Enemy_img = 4'd7;
//6'd34,6'd36,6'd62,6'd63,6'd64,6'd67,6'd68,6'd69,6'd73,6'd74,6'd75,6'd76,6'd77,6'd79,6'd82,6'd83,6'd91,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd46,6'd48,6'd96,6'd101,6'd102: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd97,6'd98,6'd99,6'd100,6'd103,6'd104,6'd105: Enemy_img = 4'd7;
//6'd36,6'd37,6'd62,6'd63,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93: Enemy_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd107: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd106: Enemy_img = 4'd7;
//6'd82,6'd84: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd60,6'd61,6'd62,6'd63,6'd64,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd78,6'd79,6'd81,6'd83,6'd85,6'd90: Enemy_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd92,6'd93,6'd95,6'd96,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd94,6'd97: Enemy_img = 4'd7;
//6'd81,6'd82,6'd83,6'd85,6'd86: Enemy_img = 4'd14;
//6'd35,6'd36,6'd39,6'd61,6'd62,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd76,6'd77,6'd84,6'd87,6'd90,6'd110,6'd111: Enemy_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92,6'd93,6'd98,6'd99,6'd104: Enemy_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd94,6'd95,6'd96,6'd97,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd7;
//6'd81,6'd82,6'd83,6'd85,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd59,6'd63,6'd66,6'd70,6'd72,6'd84,6'd86,6'd87,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd97,6'd98,6'd99: Enemy_img = 4'd6;
//6'd46,6'd49,6'd52,6'd54,6'd92,6'd93,6'd94,6'd95,6'd96,6'd100,6'd101: Enemy_img = 4'd7;
//6'd87,6'd88,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd39,6'd40,6'd41,6'd43,6'd59,6'd60,6'd61,6'd62,6'd63,6'd66,6'd67,6'd68,6'd76,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd86,6'd89,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd91,6'd97,6'd98: Enemy_img = 4'd6;
//6'd92,6'd93,6'd94,6'd95,6'd96,6'd99: Enemy_img = 4'd7;
//6'd66,6'd69,6'd76,6'd82,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd35,6'd37,6'd41,6'd44,6'd45,6'd46,6'd48,6'd51,6'd60,6'd61,6'd62,6'd63,6'd67,6'd68,6'd70,6'd71,6'd72,6'd74,6'd75,6'd77,6'd78,6'd80,6'd81,6'd89: Enemy_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd92,6'd93,6'd94,6'd95,6'd96: Enemy_img = 4'd6;
//6'd67,6'd69,6'd70,6'd71,6'd72,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85,6'd86,6'd90,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd52,6'd53,6'd57,6'd58,6'd61,6'd62,6'd63,6'd66,6'd68,6'd73,6'd74,6'd79,6'd80,6'd87,6'd88,6'd89,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd40,6'd93,6'd94: Enemy_img = 4'd6;
//6'd81: Enemy_img = 4'd9;
//6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd87,6'd88,6'd89,6'd90,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd36,6'd37,6'd47,6'd48,6'd51,6'd52,6'd56,6'd57,6'd58,6'd59,6'd63,6'd68,6'd69,6'd74,6'd75,6'd80,6'd83,6'd84,6'd85,6'd86,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43: Enemy_img = 4'd7;
//6'd81: Enemy_img = 4'd9;
//6'd82: Enemy_img = 4'd10;
//6'd69,6'd71,6'd74,6'd76,6'd77,6'd78,6'd79,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd93,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd34,6'd47,6'd50,6'd51,6'd52,6'd57,6'd58,6'd59,6'd60,6'd63,6'd65,6'd66,6'd67,6'd68,6'd70,6'd72,6'd73,6'd75,6'd84,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd39,6'd40: Enemy_img = 4'd6;
//6'd41,6'd42: Enemy_img = 4'd7;
//6'd81: Enemy_img = 4'd9;
//6'd82: Enemy_img = 4'd10;
//6'd67,6'd69,6'd77,6'd78,6'd79,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd48,6'd49,6'd51,6'd52,6'd57,6'd58,6'd61,6'd62,6'd66,6'd68,6'd70,6'd71,6'd76,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd74,6'd75: Enemy_img = 4'd2;
//6'd38,6'd39: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42: Enemy_img = 4'd7;
//6'd81,6'd82,6'd83: Enemy_img = 4'd10;
//6'd66,6'd67,6'd70,6'd71,6'd72,6'd79,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd34,6'd35,6'd47,6'd48,6'd51,6'd55,6'd56,6'd60,6'd61,6'd62,6'd65,6'd68,6'd69,6'd78,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd76,6'd77: Enemy_img = 4'd2;
//6'd40,6'd41,6'd42: Enemy_img = 4'd6;
//6'd82,6'd83: Enemy_img = 4'd9;
//6'd67,6'd71,6'd72,6'd79,6'd80,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd34,6'd35,6'd49,6'd50,6'd55,6'd56,6'd58,6'd62,6'd63,6'd64,6'd66,6'd73,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd69,6'd70,6'd77: Enemy_img = 4'd2;
//6'd42,6'd43,6'd44,6'd46: Enemy_img = 4'd6;
//6'd41: Enemy_img = 4'd7;
//6'd82: Enemy_img = 4'd9;
//6'd66,6'd75,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd34,6'd35,6'd36,6'd49,6'd50,6'd54,6'd55,6'd56,6'd58,6'd59,6'd60,6'd61,6'd63,6'd64,6'd65,6'd67,6'd74,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd76: Enemy_img = 4'd2;
//6'd45,6'd46: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43,6'd44: Enemy_img = 4'd7;
//6'd82: Enemy_img = 4'd9;
//6'd68,6'd69,6'd74,6'd78,6'd79,6'd80,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd28,6'd29,6'd35,6'd54,6'd55,6'd56,6'd59,6'd60,6'd61,6'd63,6'd65,6'd66,6'd67,6'd70,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72,6'd76: Enemy_img = 4'd2;
//6'd44,6'd45: Enemy_img = 4'd6;
//6'd40,6'd41,6'd42,6'd43: Enemy_img = 4'd7;
//6'd66,6'd67,6'd70,6'd73,6'd74,6'd78,6'd79,6'd80,6'd83,6'd84,6'd85,6'd86,6'd87,6'd88,6'd89,6'd90,6'd92,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd36,6'd37,6'd48,6'd53,6'd54,6'd57,6'd58,6'd59,6'd61,6'd65,6'd68,6'd69: Enemy_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd72: Enemy_img = 4'd2;
//6'd44,6'd45: Enemy_img = 4'd6;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd63: Enemy_img = 4'd7;
//6'd29,6'd30,6'd68,6'd69,6'd70,6'd73,6'd74,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd87,6'd88,6'd89,6'd90,6'd91,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108: Enemy_img = 4'd14;
//6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd52,6'd53,6'd55,6'd56,6'd65,6'd66,6'd67,6'd92,6'd109,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd71: Enemy_img = 4'd2;
//6'd44,6'd60,6'd61: Enemy_img = 4'd6;
//6'd41,6'd42,6'd43,6'd62: Enemy_img = 4'd7;
//6'd27,6'd28,6'd29,6'd30,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd73,6'd74,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd88,6'd89,6'd91,6'd92,6'd95,6'd96,6'd97,6'd98,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd33,6'd51,6'd54,6'd64,6'd93,6'd94,6'd100,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd43,6'd44,6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd61,6'd62,6'd63,6'd100: Enemy_img = 4'd7;
//6'd29: Enemy_img = 4'd13;
//6'd27,6'd28,6'd65,6'd66,6'd67,6'd68,6'd69,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd86,6'd88,6'd89,6'd91,6'd92,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd36,6'd37,6'd87,6'd93,6'd94,6'd95,6'd96,6'd103: Enemy_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd53,6'd55,6'd56,6'd58,6'd59,6'd60: Enemy_img = 4'd6;
//6'd57,6'd61,6'd62,6'd63,6'd64,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: Enemy_img = 4'd7;
//6'd27,6'd28: Enemy_img = 4'd13;
//6'd29,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd82,6'd83,6'd84,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd95,6'd105,6'd106,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd34,6'd36,6'd37,6'd38,6'd85,6'd86,6'd94,6'd104,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd63: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd6;
//6'd50,6'd51,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103: Enemy_img = 4'd7;
//6'd28,6'd29,6'd66,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd86,6'd87,6'd88,6'd89,6'd90,6'd91,6'd92,6'd93,6'd94,6'd107,6'd108,6'd109: Enemy_img = 4'd14;
//6'd36,6'd38,6'd39,6'd40,6'd85,6'd106,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd64: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd46,6'd55,6'd56,6'd57,6'd60: Enemy_img = 4'd6;
//6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd58,6'd59,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104: Enemy_img = 4'd7;
//6'd28,6'd29,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd79,6'd80,6'd82,6'd83,6'd84,6'd85,6'd90,6'd91,6'd92,6'd107,6'd108: Enemy_img = 4'd14;
//6'd31,6'd32,6'd34,6'd39,6'd40,6'd81,6'd86,6'd87,6'd88,6'd89,6'd106,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd65: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd45,6'd56,6'd57,6'd98,6'd99,6'd100,6'd101,6'd103,6'd106: Enemy_img = 4'd6;
//6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd58,6'd94,6'd95,6'd96,6'd97,6'd102,6'd104: Enemy_img = 4'd7;
//6'd64,6'd65,6'd68,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd87,6'd88,6'd90,6'd91,6'd92,6'd109: Enemy_img = 4'd14;
//6'd29,6'd31,6'd32,6'd34,6'd36,6'd61,6'd62,6'd63,6'd66,6'd67,6'd82,6'd86,6'd89,6'd108,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd66: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd54,6'd55,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd104,6'd105: Enemy_img = 4'd6;
//6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd93,6'd94: Enemy_img = 4'd7;
//6'd61,6'd62,6'd63,6'd67,6'd69,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd83,6'd84,6'd85,6'd87,6'd88,6'd89,6'd90: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd35,6'd36,6'd37,6'd38,6'd59,6'd60,6'd64,6'd65,6'd66,6'd82,6'd86,6'd91,6'd108,6'd109: Enemy_img = 4'd15;
//endcase
//end
//6'd67: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd44,6'd45,6'd54,6'd55,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100: Enemy_img = 4'd6;
//6'd43,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd92,6'd93,6'd94: Enemy_img = 4'd7;
//6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd77,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd86,6'd88,6'd89: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd40,6'd56,6'd57,6'd58,6'd61,6'd82,6'd83,6'd87,6'd110: Enemy_img = 4'd15;
//endcase
//end
//6'd68: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd94,6'd95,6'd96,6'd97: Enemy_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd91,6'd92,6'd93: Enemy_img = 4'd7;
//6'd57,6'd58,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd74,6'd76,6'd77,6'd78,6'd79,6'd84,6'd88,6'd89: Enemy_img = 4'd14;
//6'd30,6'd31,6'd32,6'd35,6'd36,6'd39,6'd40,6'd59,6'd60,6'd61,6'd69,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd69: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd41,6'd42,6'd43,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd35,6'd36,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd91,6'd92: Enemy_img = 4'd7;
//6'd57,6'd59,6'd60,6'd65,6'd66,6'd67,6'd70,6'd71,6'd72,6'd73,6'd76,6'd77,6'd80,6'd81,6'd82,6'd86,6'd87,6'd88,6'd89: Enemy_img = 4'd14;
//6'd28,6'd30,6'd31,6'd32,6'd33,6'd54,6'd55,6'd56,6'd58,6'd61,6'd62,6'd63,6'd64,6'd69,6'd78,6'd79,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd70: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd39,6'd41,6'd42,6'd45,6'd46,6'd47,6'd92,6'd93,6'd94,6'd95: Enemy_img = 4'd6;
//6'd35,6'd36,6'd37,6'd40,6'd43,6'd44,6'd48,6'd49,6'd90,6'd91: Enemy_img = 4'd7;
//6'd56,6'd58,6'd60,6'd62,6'd63,6'd72,6'd73,6'd74,6'd75,6'd76,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd28,6'd29,6'd31,6'd32,6'd33,6'd52,6'd53,6'd54,6'd55,6'd57,6'd59,6'd61,6'd64,6'd65,6'd66,6'd69,6'd70,6'd71,6'd77,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd71: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd46,6'd47,6'd48,6'd92,6'd93,6'd94: Enemy_img = 4'd6;
//6'd39,6'd45,6'd90,6'd91: Enemy_img = 4'd7;
//6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd70,6'd72,6'd74,6'd75,6'd76,6'd77,6'd79,6'd80,6'd81,6'd82,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd51,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd69,6'd71,6'd73,6'd78,6'd83,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd72: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd37,6'd38,6'd49,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd35,6'd48,6'd90: Enemy_img = 4'd7;
//6'd42,6'd64,6'd65,6'd66,6'd67,6'd69,6'd70,6'd73,6'd75,6'd78,6'd79,6'd80,6'd84,6'd86: Enemy_img = 4'd14;
//6'd27,6'd29,6'd31,6'd32,6'd43,6'd44,6'd45,6'd52,6'd61,6'd62,6'd63,6'd68,6'd71,6'd72,6'd74,6'd76,6'd77,6'd81,6'd82,6'd83,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd73: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd48,6'd49,6'd91,6'd92,6'd93: Enemy_img = 4'd6;
//6'd35,6'd37,6'd38,6'd89,6'd90: Enemy_img = 4'd7;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd55,6'd67,6'd70,6'd72,6'd73,6'd77,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84: Enemy_img = 4'd14;
//6'd26,6'd28,6'd30,6'd31,6'd32,6'd33,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd56,6'd57,6'd58,6'd59,6'd60,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd71,6'd74,6'd75,6'd76,6'd81,6'd85,6'd87,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd74: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd34,6'd35,6'd36,6'd49,6'd50,6'd91,6'd92: Enemy_img = 4'd6;
//6'd37,6'd38,6'd90: Enemy_img = 4'd7;
//6'd32,6'd33,6'd40,6'd41,6'd42,6'd56,6'd57,6'd59,6'd60,6'd61,6'd70,6'd72,6'd73,6'd75,6'd78,6'd79,6'd80,6'd82,6'd83,6'd84,6'd88: Enemy_img = 4'd14;
//6'd26,6'd29,6'd30,6'd31,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55,6'd58,6'd62,6'd63,6'd65,6'd66,6'd67,6'd77,6'd81,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd75: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd36,6'd49,6'd50,6'd51,6'd90,6'd91: Enemy_img = 4'd6;
//6'd37,6'd89: Enemy_img = 4'd7;
//6'd31,6'd32,6'd33,6'd39,6'd40,6'd41,6'd45,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd87,6'd88: Enemy_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd44,6'd46,6'd47,6'd54,6'd55,6'd56,6'd57,6'd64,6'd68,6'd69,6'd70,6'd71,6'd72,6'd74,6'd76,6'd81,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd76: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd54,6'd90,6'd91: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd66,6'd67,6'd89: Enemy_img = 4'd7;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd41,6'd42,6'd44,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd74,6'd77,6'd79,6'd86,6'd87: Enemy_img = 4'd14;
//6'd24,6'd25,6'd26,6'd43,6'd45,6'd46,6'd47,6'd56,6'd65,6'd70,6'd71,6'd72,6'd73,6'd75,6'd76,6'd78,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd77: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd90,6'd91: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd66,6'd67,6'd68,6'd69: Enemy_img = 4'd7;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd83,6'd85,6'd87,6'd88: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd47,6'd55,6'd73,6'd74,6'd75,6'd84,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd78: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd89,6'd90: Enemy_img = 4'd6;
//6'd48,6'd49,6'd50,6'd51,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72: Enemy_img = 4'd7;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd78,6'd79,6'd80,6'd81,6'd84,6'd85,6'd87: Enemy_img = 4'd14;
//6'd22,6'd23,6'd25,6'd46,6'd55,6'd75,6'd76,6'd77,6'd82,6'd83,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd79: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd52,6'd53,6'd90: Enemy_img = 4'd6;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd75: Enemy_img = 4'd7;
//6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd43,6'd44,6'd57,6'd58,6'd59,6'd60,6'd82,6'd84,6'd85,6'd87: Enemy_img = 4'd14;
//6'd28,6'd29,6'd30,6'd33,6'd42,6'd45,6'd54,6'd55,6'd56,6'd78,6'd79,6'd80,6'd81,6'd83,6'd86,6'd88: Enemy_img = 4'd15;
//endcase
//end
//6'd80: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd89: Enemy_img = 4'd6;
//6'd50,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77: Enemy_img = 4'd7;
//6'd35,6'd36,6'd37,6'd39,6'd40,6'd43,6'd44,6'd59,6'd60,6'd61,6'd81,6'd82,6'd83: Enemy_img = 4'd14;
//6'd32,6'd33,6'd34,6'd38,6'd41,6'd42,6'd45,6'd46,6'd47,6'd55,6'd56,6'd57,6'd58,6'd79,6'd80,6'd84,6'd85,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd81: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd52,6'd72,6'd89: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78: Enemy_img = 4'd7;
//6'd37,6'd42,6'd44,6'd45,6'd46,6'd58,6'd82,6'd83,6'd86,6'd87: Enemy_img = 4'd14;
//6'd35,6'd36,6'd38,6'd39,6'd41,6'd43,6'd47,6'd48,6'd49,6'd57,6'd59,6'd81,6'd84,6'd85: Enemy_img = 4'd15;
//endcase
//end
//6'd82: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd51,6'd67,6'd68,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd89: Enemy_img = 4'd6;
//6'd52,6'd53,6'd54,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd69,6'd77,6'd78,6'd79: Enemy_img = 4'd7;
//6'd41,6'd42,6'd46,6'd47,6'd48,6'd83,6'd84,6'd87: Enemy_img = 4'd14;
//6'd36,6'd38,6'd40,6'd43,6'd44,6'd45,6'd49,6'd56,6'd57,6'd58,6'd81,6'd82,6'd85,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd83: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd50,6'd51,6'd52,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd81: Enemy_img = 4'd6;
//6'd53,6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd7;
//6'd43,6'd44,6'd45,6'd47,6'd57,6'd58,6'd59,6'd85: Enemy_img = 4'd14;
//6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd46,6'd48,6'd56,6'd84,6'd86,6'd87: Enemy_img = 4'd15;
//endcase
//end
//6'd84: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd53,6'd54,6'd65,6'd66,6'd67,6'd68,6'd69,6'd70,6'd71,6'd72,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd7;
//6'd36,6'd37,6'd38,6'd39,6'd45,6'd57,6'd58,6'd85,6'd86,6'd87: Enemy_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd46,6'd47,6'd48,6'd49,6'd50,6'd55,6'd56,6'd84: Enemy_img = 4'd15;
//endcase
//end
//6'd85: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd69,6'd80,6'd82,6'd84: Enemy_img = 4'd6;
//6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd39,6'd40: Enemy_img = 4'd13;
//6'd37,6'd38,6'd47,6'd48,6'd57,6'd58,6'd87,6'd88: Enemy_img = 4'd14;
//6'd43,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd55,6'd56,6'd86: Enemy_img = 4'd15;
//endcase
//end
//6'd86: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd63,6'd64,6'd65,6'd66,6'd67: Enemy_img = 4'd6;
//6'd59,6'd60,6'd61,6'd62: Enemy_img = 4'd7;
//6'd37,6'd38: Enemy_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd47,6'd48,6'd49,6'd50,6'd56,6'd87: Enemy_img = 4'd14;
//6'd44,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57: Enemy_img = 4'd15;
//endcase
//end
//6'd87: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd62,6'd63,6'd64,6'd65: Enemy_img = 4'd6;
//6'd58,6'd59,6'd60,6'd61: Enemy_img = 4'd7;
//6'd38,6'd39,6'd40,6'd41,6'd49,6'd50,6'd51,6'd53,6'd55,6'd56,6'd57,6'd88: Enemy_img = 4'd14;
//6'd46,6'd47,6'd48,6'd52,6'd54: Enemy_img = 4'd15;
//endcase
//end
//6'd88: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd61,6'd62,6'd63,6'd64: Enemy_img = 4'd6;
//6'd59,6'd60: Enemy_img = 4'd7;
//6'd38,6'd39,6'd49,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd40,6'd41,6'd47,6'd48,6'd50: Enemy_img = 4'd15;
//endcase
//end
//6'd89: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61,6'd62: Enemy_img = 4'd6;
//6'd58,6'd59: Enemy_img = 4'd7;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd39,6'd48,6'd49: Enemy_img = 4'd15;
//endcase
//end
//6'd90: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd60,6'd61: Enemy_img = 4'd6;
//6'd58,6'd59: Enemy_img = 4'd7;
//6'd52,6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd50,6'd51,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd91: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd59,6'd60: Enemy_img = 4'd6;
//6'd53,6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd50,6'd51,6'd52: Enemy_img = 4'd15;
//endcase
//end
//6'd92: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58,6'd59: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56: Enemy_img = 4'd14;
//6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd93: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57: Enemy_img = 4'd14;
//6'd52,6'd53: Enemy_img = 4'd15;
//endcase
//end
//6'd94: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd58: Enemy_img = 4'd6;
//6'd54,6'd55,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd95: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd55: Enemy_img = 4'd14;
//6'd54,6'd56: Enemy_img = 4'd15;
//endcase
//end
//6'd96: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd97: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd98: begin
//case(x)
//default: Enemy_img = 4'd0;
//6'd56: Enemy_img = 4'd14;
//endcase
//end
//6'd99: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd100: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd101: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd102: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd103: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd104: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd105: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd106: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd107: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd108: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd109: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd110: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd111: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd112: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd113: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd114: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd115: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd116: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd117: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd118: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd119: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd120: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd121: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd122: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd123: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd124: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd125: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd126: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//6'd127: begin
//case(x)
//default: Enemy_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//
//endcase


end
endfunction
function [3:0] Bullet_img(input [6:0] x, input [6:0] y, input [3:0] angle, input [1:0] b_type);
begin

//case(b_type)
//
//2'd0: begin
//case(angle)
//// Bullet_type_0 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd9,6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd2;
//6'd8,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd18,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd0;
//default: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd2;
//6'd9: Bullet_img = 4'd3;
//6'd8,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd1;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd19: Bullet_img = 4'd1;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd20,6'd21: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd24: Bullet_img = 4'd4;
//6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd13,6'd14,6'd15,6'd16,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd1;
//6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd18: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd1;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd19: Bullet_img = 4'd1;
//6'd7,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd20,6'd21: Bullet_img = 4'd4;
//6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd19: Bullet_img = 4'd1;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13: Bullet_img = 4'd1;
//6'd9: Bullet_img = 4'd3;
//6'd8,6'd10,6'd11,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11: Bullet_img = 4'd1;
//6'd8,6'd12,6'd13,6'd14: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd1;
//6'd11: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd1;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd1;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd21: Bullet_img = 4'd3;
//6'd18,6'd19,6'd22: Bullet_img = 4'd4;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd21: Bullet_img = 4'd3;
//6'd17,6'd18,6'd20,6'd22,6'd23: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd22: Bullet_img = 4'd2;
//6'd16,6'd17,6'd19,6'd20,6'd21,6'd24: Bullet_img = 4'd4;
//6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd4;
//6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd14,6'd15,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd14: Bullet_img = 4'd2;
//6'd11,6'd12,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd13,6'd14: Bullet_img = 4'd2;
//6'd11,6'd15,6'd17,6'd18: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd1;
//6'd12,6'd13: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd1;
//6'd11,6'd12: Bullet_img = 4'd2;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11: Bullet_img = 4'd2;
//6'd12,6'd14,6'd15: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd2;
//6'd11: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd20: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd3;
//6'd16,6'd19,6'd21,6'd22: Bullet_img = 4'd4;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd20: Bullet_img = 4'd2;
//6'd16,6'd18,6'd19: Bullet_img = 4'd4;
//6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd15,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd15,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd14,6'd15,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14: Bullet_img = 4'd1;
//6'd15: Bullet_img = 4'd2;
//6'd12: Bullet_img = 4'd4;
//6'd16,6'd17,6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd14: Bullet_img = 4'd2;
//6'd12,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd14: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd13: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd13: Bullet_img = 4'd2;
//6'd14: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd13: Bullet_img = 4'd2;
//6'd14: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd2;
//6'd13: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15: Bullet_img = 4'd1;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd3;
//6'd17: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15: Bullet_img = 4'd1;
//6'd16: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd16: Bullet_img = 4'd2;
//6'd14,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd16: Bullet_img = 4'd2;
//6'd14,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd16: Bullet_img = 4'd2;
//6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd16: Bullet_img = 4'd2;
//6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd16: Bullet_img = 4'd2;
//6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd2;
//6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd4;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12: Bullet_img = 4'd1;
//6'd13: Bullet_img = 4'd3;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd11,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd12,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd12,6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd12,6'd13,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd13,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd13,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14,6'd16,6'd19: Bullet_img = 4'd4;
//6'd17,6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//6'd14,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd15,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd17,6'd18: Bullet_img = 4'd2;
//6'd15,6'd19: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd19: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd19: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd13;
//6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd2;
//6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd4;
//6'd12,6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd2;
//6'd10,6'd11,6'd13,6'd14: Bullet_img = 4'd4;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd1;
//6'd10: Bullet_img = 4'd3;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd10: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd1;
//6'd10,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd10,6'd11,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd11,6'd12,6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd12,6'd13,6'd15,6'd16,6'd17,6'd19,6'd20: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd13,6'd14,6'd16,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd2;
//6'd14,6'd15,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd1;
//6'd18,6'd19: Bullet_img = 4'd2;
//6'd20: Bullet_img = 4'd4;
//6'd21: Bullet_img = 4'd13;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd18: Bullet_img = 4'd1;
//6'd19,6'd20: Bullet_img = 4'd2;
//6'd17,6'd21: Bullet_img = 4'd4;
//6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd20,6'd21: Bullet_img = 4'd2;
//6'd17,6'd18,6'd22: Bullet_img = 4'd4;
//6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd21,6'd22: Bullet_img = 4'd2;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd2;
//6'd9,6'd11,6'd12,6'd13: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9: Bullet_img = 4'd1;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd11: Bullet_img = 4'd1;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd19,6'd20: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14: Bullet_img = 4'd1;
//6'd10,6'd11,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd12,6'd13,6'd14,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd22,6'd23: Bullet_img = 4'd13;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd15,6'd16,6'd22,6'd23: Bullet_img = 4'd4;
//6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd20,6'd21: Bullet_img = 4'd1;
//6'd22,6'd23: Bullet_img = 4'd2;
//6'd19,6'd24: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd1;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd2;
//6'd21: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd17,6'd18,6'd20: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd1;
//6'd20,6'd21: Bullet_img = 4'd2;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd1;
//6'd19,6'd20: Bullet_img = 4'd2;
//6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd18,6'd19: Bullet_img = 4'd2;
//6'd14,6'd15,6'd17,6'd21: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd13,6'd14,6'd15,6'd16,6'd20,6'd21: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd1;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd18: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd16,6'd17: Bullet_img = 4'd4;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd10: Bullet_img = 4'd2;
//6'd8,6'd11,6'd12,6'd13,6'd15,6'd16: Bullet_img = 4'd4;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd11: Bullet_img = 4'd3;
//6'd9,6'd10,6'd12,6'd14,6'd15: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd11: Bullet_img = 4'd3;
//6'd10,6'd13,6'd14: Bullet_img = 4'd4;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd1;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd2;
//6'd19: Bullet_img = 4'd4;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd18: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16,6'd17,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd20: Bullet_img = 4'd4;
//6'd14,6'd15,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd13,6'd14,6'd15,6'd16,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd12,6'd13,6'd14,6'd15,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd12,6'd13,6'd14,6'd15,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd12: Bullet_img = 4'd2;
//6'd13,6'd14,6'd16: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd12: Bullet_img = 4'd2;
//6'd14: Bullet_img = 4'd3;
//6'd10,6'd11,6'd13,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd1;
//6'd12,6'd13: Bullet_img = 4'd4;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19: Bullet_img = 4'd1;
//6'd17: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd15: Bullet_img = 4'd2;
//6'd17: Bullet_img = 4'd3;
//6'd16: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd2;
//6'd12: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14: Bullet_img = 4'd2;
//6'd13: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd13;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd1;
//6'd14: Bullet_img = 4'd2;
//6'd13: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd14,6'd15: Bullet_img = 4'd2;
//6'd13,6'd17: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd15: Bullet_img = 4'd2;
//6'd13,6'd14,6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18: Bullet_img = 4'd1;
//6'd15: Bullet_img = 4'd2;
//6'd12,6'd13,6'd14: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd4;
//6'd16,6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd13,6'd16,6'd18: Bullet_img = 4'd4;
//6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd21: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd3;
//6'd16,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd10,6'd11: Bullet_img = 4'd2;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd1;
//6'd11,6'd12: Bullet_img = 4'd2;
//6'd10,6'd14,6'd15: Bullet_img = 4'd4;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd16: Bullet_img = 4'd1;
//6'd12,6'd13: Bullet_img = 4'd2;
//6'd11,6'd15: Bullet_img = 4'd4;
//6'd10: Bullet_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd1;
//6'd13,6'd14: Bullet_img = 4'd2;
//6'd12: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd13;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd17,6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd14,6'd16,6'd18,6'd19: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd12,6'd13,6'd15,6'd16,6'd17,6'd19,6'd20: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd20,6'd21: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd21,6'd22: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd22: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd24: Bullet_img = 4'd1;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd1;
//6'd21,6'd22: Bullet_img = 4'd3;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd2;
//6'd18,6'd19,6'd21,6'd22: Bullet_img = 4'd4;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd4;
//6'd19,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd4;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11: Bullet_img = 4'd1;
//6'd8: Bullet_img = 4'd2;
//6'd13,6'd14: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd1;
//6'd9,6'd10,6'd11: Bullet_img = 4'd2;
//6'd8: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd16: Bullet_img = 4'd1;
//6'd12,6'd13: Bullet_img = 4'd2;
//6'd9,6'd10,6'd11,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd1;
//6'd14: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd16,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd9,6'd10: Bullet_img = 4'd13;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd15,6'd16,6'd17,6'd18,6'd22,6'd23: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd25: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd1;
//6'd23: Bullet_img = 4'd3;
//6'd13,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd4;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd2;
//6'd18,6'd19,6'd20,6'd21,6'd24: Bullet_img = 4'd4;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd23: Bullet_img = 4'd4;
//6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd4;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd25: Bullet_img = 4'd1;
//6'd12,6'd13,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd1;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//6'd24: Bullet_img = 4'd3;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd0;
//default: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd2;
//6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25: Bullet_img = 4'd4;
//6'd9,6'd10,6'd11: Bullet_img = 4'd13;
//6'd8,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25: Bullet_img = 4'd4;
//6'd15,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_0 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd1;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd1;
//6'd21: Bullet_img = 4'd4;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23: Bullet_img = 4'd1;
//6'd18,6'd19,6'd20,6'd24: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd1;
//6'd23: Bullet_img = 4'd3;
//6'd16,6'd17,6'd18,6'd21,6'd22,6'd24: Bullet_img = 4'd4;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd16,6'd17,6'd18: Bullet_img = 4'd1;
//6'd15,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd15: Bullet_img = 4'd1;
//6'd11,6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25: Bullet_img = 4'd4;
//6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd14,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11: Bullet_img = 4'd2;
//6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8: Bullet_img = 4'd2;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd13,6'd14: Bullet_img = 4'd4;
//6'd9,6'd10,6'd11: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//2'd1: begin
//case(angle)
//// Bullet_type_1 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd2;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd1;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11: Bullet_img = 4'd2;
//6'd8,6'd9: Bullet_img = 4'd3;
//6'd43: Bullet_img = 4'd13;
//6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd14,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd2;
//6'd7,6'd8,6'd10: Bullet_img = 4'd3;
//6'd9: Bullet_img = 4'd4;
//default: Bullet_img = 4'd12;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd14,6'd44,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd6,6'd43: Bullet_img = 4'd1;
//6'd11,6'd12,6'd13,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd2;
//6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd3;
//default: Bullet_img = 4'd12;
//6'd4,6'd5,6'd45: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd14,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd12,6'd13,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44: Bullet_img = 4'd2;
//6'd6,6'd8,6'd9,6'd10,6'd11,6'd43: Bullet_img = 4'd3;
//6'd7,6'd25: Bullet_img = 4'd4;
//default: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd14,6'd43,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd2;
//6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd3;
//6'd44: Bullet_img = 4'd8;
//6'd26: Bullet_img = 4'd12;
//default: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11: Bullet_img = 4'd2;
//6'd8,6'd9: Bullet_img = 4'd3;
//6'd43: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11: Bullet_img = 4'd2;
//6'd8,6'd9: Bullet_img = 4'd3;
//6'd43: Bullet_img = 4'd13;
//6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd2;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd2;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd1;
//6'd39,6'd40: Bullet_img = 4'd2;
//6'd43: Bullet_img = 4'd13;
//6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd42: Bullet_img = 4'd2;
//6'd41: Bullet_img = 4'd3;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd2;
//6'd41: Bullet_img = 4'd3;
//6'd43: Bullet_img = 4'd8;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd2;
//6'd31,6'd32: Bullet_img = 4'd12;
//6'd42: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd12;
//6'd42: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd12;
//6'd32,6'd33: Bullet_img = 4'd13;
//6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd34: Bullet_img = 4'd2;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd2;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd2;
//6'd25: Bullet_img = 4'd4;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd26: Bullet_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd1;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd12;
//6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd9: Bullet_img = 4'd3;
//6'd15,6'd16: Bullet_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd8,6'd9,6'd10: Bullet_img = 4'd3;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//6'd7,6'd8,6'd10: Bullet_img = 4'd3;
//6'd9: Bullet_img = 4'd4;
//6'd16,6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7: Bullet_img = 4'd1;
//6'd13,6'd14,6'd20,6'd21: Bullet_img = 4'd2;
//6'd8,6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd3;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7: Bullet_img = 4'd1;
//6'd12,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//6'd8: Bullet_img = 4'd4;
//6'd5,6'd6: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd7,6'd8,6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd10,6'd11: Bullet_img = 4'd3;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd2;
//6'd10: Bullet_img = 4'd3;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34: Bullet_img = 4'd3;
//6'd39: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd2;
//6'd33,6'd34,6'd35,6'd37: Bullet_img = 4'd3;
//6'd36: Bullet_img = 4'd4;
//6'd38: Bullet_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd3;
//6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd32: Bullet_img = 4'd2;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd3;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd32: Bullet_img = 4'd2;
//6'd33,6'd34,6'd35,6'd37,6'd38: Bullet_img = 4'd3;
//6'd36: Bullet_img = 4'd4;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd36: Bullet_img = 4'd2;
//6'd35,6'd37: Bullet_img = 4'd3;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36: Bullet_img = 4'd1;
//6'd25,6'd33: Bullet_img = 4'd2;
//6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32: Bullet_img = 4'd12;
//6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//6'd28,6'd29: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd2;
//6'd23: Bullet_img = 4'd4;
//6'd22,6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd12;
//6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd12;
//6'd16,6'd17,6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd2;
//6'd18,6'd19: Bullet_img = 4'd12;
//6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd12;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd2;
//6'd9: Bullet_img = 4'd13;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd12,6'd13: Bullet_img = 4'd2;
//6'd11: Bullet_img = 4'd3;
//6'd9: Bullet_img = 4'd8;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd13: Bullet_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd1;
//6'd27,6'd29,6'd30,6'd31: Bullet_img = 4'd3;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd31,6'd32: Bullet_img = 4'd3;
//6'd30: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26: Bullet_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd3;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd2;
//6'd28,6'd29,6'd30,6'd32,6'd33: Bullet_img = 4'd3;
//6'd31: Bullet_img = 4'd4;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd2;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd3;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd1;
//6'd20,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd29,6'd30: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd28: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd28,6'd29: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd27,6'd28,6'd29: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd4;
//6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd24,6'd25: Bullet_img = 4'd12;
//6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd19,6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd2;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//6'd20,6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//6'd14,6'd15: Bullet_img = 4'd13;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd3;
//6'd15: Bullet_img = 4'd8;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd2;
//6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd1;
//6'd24: Bullet_img = 4'd3;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd25,6'd26: Bullet_img = 4'd3;
//6'd24: Bullet_img = 4'd4;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd3;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd27: Bullet_img = 4'd3;
//6'd26: Bullet_img = 4'd4;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd27: Bullet_img = 4'd2;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd3;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28: Bullet_img = 4'd1;
//6'd21,6'd22,6'd23,6'd25,6'd26,6'd27: Bullet_img = 4'd2;
//6'd24: Bullet_img = 4'd3;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd4;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd25,6'd26: Bullet_img = 4'd12;
//6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//6'd21,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd1;
//6'd24: Bullet_img = 4'd3;
//6'd21,6'd22,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd2;
//6'd23: Bullet_img = 4'd8;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd1;
//6'd16,6'd19: Bullet_img = 4'd3;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd18,6'd19,6'd20: Bullet_img = 4'd3;
//6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd20,6'd21: Bullet_img = 4'd3;
//6'd19: Bullet_img = 4'd4;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd1;
//6'd21: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd3;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd3;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd3;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd25,6'd26,6'd27: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd19,6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27: Bullet_img = 4'd2;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd25: Bullet_img = 4'd2;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd20,6'd21: Bullet_img = 4'd13;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd4;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd25,6'd26: Bullet_img = 4'd12;
//6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29: Bullet_img = 4'd2;
//6'd28: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd33: Bullet_img = 4'd13;
//6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd1;
//6'd29: Bullet_img = 4'd2;
//6'd30,6'd31: Bullet_img = 4'd3;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd2;
//6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30: Bullet_img = 4'd8;
//6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd3;
//6'd10,6'd11: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd1;
//6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd3;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd1;
//6'd15,6'd16: Bullet_img = 4'd2;
//6'd12,6'd13: Bullet_img = 4'd3;
//6'd11,6'd14: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd3;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd22,6'd23: Bullet_img = 4'd2;
//6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd3;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd15,6'd16,6'd17,6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd10,6'd11,6'd13,6'd14: Bullet_img = 4'd3;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd12;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd15,6'd22,6'd23: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19: Bullet_img = 4'd12;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20: Bullet_img = 4'd12;
//6'd16,6'd17: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd12;
//6'd17,6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22: Bullet_img = 4'd12;
//6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd2;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd16: Bullet_img = 4'd2;
//6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//6'd12: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd4;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd23,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd27,6'd28: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32: Bullet_img = 4'd12;
//6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd2;
//6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd39: Bullet_img = 4'd13;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd2;
//6'd37: Bullet_img = 4'd3;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd2;
//6'd39: Bullet_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37: Bullet_img = 4'd8;
//6'd35: Bullet_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7,6'd13: Bullet_img = 4'd1;
//6'd12,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//6'd5,6'd6: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd7,6'd8,6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//6'd7,6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//6'd8: Bullet_img = 4'd4;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//6'd8,6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//6'd16,6'd17: Bullet_img = 4'd12;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13: Bullet_img = 4'd2;
//6'd8,6'd9,6'd10,6'd11: Bullet_img = 4'd3;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd12;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd8,6'd9: Bullet_img = 4'd3;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd12;
//6'd15,6'd16: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10: Bullet_img = 4'd2;
//6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd12;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd34: Bullet_img = 4'd2;
//6'd25,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd12;
//6'd24,6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd32,6'd33: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd13;
//6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd2;
//6'd31,6'd32,6'd42: Bullet_img = 4'd13;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd2;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd1;
//6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd2;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39: Bullet_img = 4'd2;
//6'd41: Bullet_img = 4'd3;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd8;
//6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd13;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd38: Bullet_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38: Bullet_img = 4'd2;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd38: Bullet_img = 4'd2;
//6'd37: Bullet_img = 4'd3;
//6'd39: Bullet_img = 4'd8;
//6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd39: Bullet_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd2;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd30: Bullet_img = 4'd12;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//6'd29,6'd30: Bullet_img = 4'd12;
//6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd12;
//6'd30,6'd31,6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd2;
//6'd25: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24,6'd26: Bullet_img = 4'd12;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd2;
//6'd19,6'd20: Bullet_img = 4'd12;
//6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19: Bullet_img = 4'd12;
//6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd12;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd1;
//6'd15,6'd23: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd22,6'd23,6'd24: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd14,6'd15,6'd16,6'd17,6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd11,6'd13: Bullet_img = 4'd3;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd22,6'd23,6'd24: Bullet_img = 4'd2;
//6'd10,6'd11,6'd13,6'd14,6'd15: Bullet_img = 4'd3;
//6'd12: Bullet_img = 4'd4;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd23,6'd24: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd3;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd3;
//6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd2;
//6'd11,6'd13,6'd14,6'd15: Bullet_img = 4'd3;
//6'd12: Bullet_img = 4'd4;
//6'd10: Bullet_img = 4'd13;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15: Bullet_img = 4'd3;
//6'd9: Bullet_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd2;
//6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd1;
//6'd29: Bullet_img = 4'd2;
//6'd32: Bullet_img = 4'd3;
//6'd33: Bullet_img = 4'd8;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd33,6'd34: Bullet_img = 4'd13;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd26: Bullet_img = 4'd12;
//6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd24,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd2;
//6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd2;
//6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd2;
//6'd19,6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd2;
//6'd19,6'd20: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27: Bullet_img = 4'd2;
//6'd20: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd2;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd18,6'd19,6'd20,6'd21,6'd28: Bullet_img = 4'd2;
//6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd2;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd3;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd15,6'd16,6'd18,6'd19,6'd20: Bullet_img = 4'd3;
//6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd2;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd3;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd19,6'd20,6'd21: Bullet_img = 4'd3;
//6'd18: Bullet_img = 4'd4;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd17,6'd18,6'd19,6'd21: Bullet_img = 4'd3;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd2;
//6'd26: Bullet_img = 4'd8;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd1;
//6'd25: Bullet_img = 4'd3;
//6'd22,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//6'd22,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd26: Bullet_img = 4'd12;
//6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd4;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21,6'd29,6'd30: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21,6'd29,6'd30: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd2;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd1;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd28: Bullet_img = 4'd2;
//6'd25: Bullet_img = 4'd3;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd27,6'd28: Bullet_img = 4'd2;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd3;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd3;
//6'd23: Bullet_img = 4'd4;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd3;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd26: Bullet_img = 4'd3;
//6'd25: Bullet_img = 4'd4;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd1;
//6'd25: Bullet_img = 4'd3;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd8;
//6'd16: Bullet_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd2;
//6'd19,6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd2;
//6'd17,6'd18: Bullet_img = 4'd3;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//6'd15: Bullet_img = 4'd13;
//6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd2;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd2;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd2;
//6'd20: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd12;
//6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd23,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd25: Bullet_img = 4'd12;
//6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd4;
//6'd22,6'd23: Bullet_img = 4'd12;
//6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd2;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28: Bullet_img = 4'd13;
//6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd29,6'd30: Bullet_img = 4'd2;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd32: Bullet_img = 4'd2;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//6'd30: Bullet_img = 4'd3;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29: Bullet_img = 4'd2;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd3;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26: Bullet_img = 4'd1;
//6'd27: Bullet_img = 4'd2;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd3;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd30,6'd31,6'd32: Bullet_img = 4'd3;
//6'd29: Bullet_img = 4'd4;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd32: Bullet_img = 4'd3;
//6'd31: Bullet_img = 4'd4;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd1;
//6'd29,6'd32: Bullet_img = 4'd3;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd8;
//6'd13: Bullet_img = 4'd13;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11: Bullet_img = 4'd2;
//6'd9: Bullet_img = 4'd13;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13: Bullet_img = 4'd2;
//6'd11: Bullet_img = 4'd3;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd2;
//6'd9: Bullet_img = 4'd13;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd2;
//6'd18: Bullet_img = 4'd13;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd12;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19: Bullet_img = 4'd12;
//6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd12;
//6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd24: Bullet_img = 4'd12;
//6'd22,6'd23: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd4;
//6'd21,6'd22: Bullet_img = 4'd12;
//6'd23,6'd25: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd34,6'd35: Bullet_img = 4'd2;
//6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26: Bullet_img = 4'd13;
//6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd2;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33: Bullet_img = 4'd2;
//6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd12;
//6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd12;
//6'd30,6'd31,6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd33,6'd36: Bullet_img = 4'd2;
//6'd29,6'd30: Bullet_img = 4'd12;
//6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd30: Bullet_img = 4'd12;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd36: Bullet_img = 4'd2;
//6'd34,6'd35,6'd37,6'd38: Bullet_img = 4'd3;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd32,6'd33: Bullet_img = 4'd2;
//6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd3;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd2;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd3;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd1;
//6'd32,6'd33: Bullet_img = 4'd2;
//6'd35,6'd36: Bullet_img = 4'd3;
//6'd34,6'd37: Bullet_img = 4'd4;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd3;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34: Bullet_img = 4'd3;
//6'd37: Bullet_img = 4'd13;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38: Bullet_img = 4'd13;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8: Bullet_img = 4'd13;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7: Bullet_img = 4'd8;
//6'd8: Bullet_img = 4'd13;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd6,6'd8,6'd9: Bullet_img = 4'd2;
//6'd7: Bullet_img = 4'd3;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7: Bullet_img = 4'd1;
//6'd8,6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd2;
//6'd5: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7: Bullet_img = 4'd1;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd2;
//6'd6,6'd16,6'd17: Bullet_img = 4'd13;
//6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd34,6'd35: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd15,6'd16: Bullet_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd23: Bullet_img = 4'd12;
//6'd20,6'd21,6'd22,6'd24: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34: Bullet_img = 4'd2;
//6'd24: Bullet_img = 4'd4;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd12;
//6'd22,6'd23,6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd2;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd39,6'd40,6'd41: Bullet_img = 4'd3;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd12;
//6'd32,6'd33: Bullet_img = 4'd13;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd38,6'd39,6'd40: Bullet_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd12;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd3;
//6'd31,6'd32: Bullet_img = 4'd12;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39,6'd41: Bullet_img = 4'd3;
//6'd40: Bullet_img = 4'd4;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd36: Bullet_img = 4'd2;
//6'd37,6'd39,6'd40,6'd41: Bullet_img = 4'd3;
//6'd38: Bullet_img = 4'd4;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd41: Bullet_img = 4'd1;
//6'd28,6'd29,6'd30,6'd36: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd3;
//6'd42,6'd43: Bullet_img = 4'd13;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//6'd38: Bullet_img = 4'd3;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd2;
//6'd40,6'd41: Bullet_img = 4'd3;
//6'd6: Bullet_img = 4'd13;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd2;
//6'd40,6'd41: Bullet_img = 4'd3;
//6'd6: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd6,6'd35,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd3;
//6'd5: Bullet_img = 4'd8;
//6'd23: Bullet_img = 4'd12;
//default: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd35,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd5,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd36,6'd37: Bullet_img = 4'd2;
//6'd6,6'd38,6'd39,6'd40,6'd41,6'd43: Bullet_img = 4'd3;
//6'd24,6'd42: Bullet_img = 4'd4;
//default: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd5,6'd35,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd6,6'd43: Bullet_img = 4'd1;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd3;
//default: Bullet_img = 4'd12;
//6'd4,6'd44,6'd45: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd35,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd39,6'd41,6'd42: Bullet_img = 4'd3;
//6'd40: Bullet_img = 4'd4;
//default: Bullet_img = 4'd12;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd2;
//6'd40,6'd41: Bullet_img = 4'd3;
//6'd6: Bullet_img = 4'd13;
//6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38: Bullet_img = 4'd1;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_1 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd2;
//6'd38: Bullet_img = 4'd3;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd36: Bullet_img = 4'd2;
//6'd37,6'd38: Bullet_img = 4'd3;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd35,6'd36: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd3;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd1;
//6'd27,6'd28,6'd29,6'd30,6'd36: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39: Bullet_img = 4'd3;
//6'd40: Bullet_img = 4'd4;
//6'd42,6'd43: Bullet_img = 4'd13;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd1;
//6'd27,6'd28,6'd34,6'd35: Bullet_img = 4'd2;
//6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd3;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd38,6'd40,6'd41: Bullet_img = 4'd3;
//6'd39: Bullet_img = 4'd4;
//6'd31,6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd38,6'd39,6'd40: Bullet_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd13;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd2;
//6'd39: Bullet_img = 4'd3;
//6'd32,6'd33: Bullet_img = 4'd12;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38: Bullet_img = 4'd1;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd12;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd2;
//6'd23: Bullet_img = 4'd4;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd12;
//6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd12;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd12;
//6'd15,6'd16: Bullet_img = 4'd13;
//6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd12;
//6'd6: Bullet_img = 4'd13;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd2;
//6'd16,6'd17: Bullet_img = 4'd12;
//6'd6: Bullet_img = 4'd13;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//6'd7: Bullet_img = 4'd3;
//6'd5: Bullet_img = 4'd8;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd6,6'd8,6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd2;
//6'd7: Bullet_img = 4'd3;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7: Bullet_img = 4'd1;
//6'd8,6'd9: Bullet_img = 4'd2;
//6'd5: Bullet_img = 4'd13;
//6'd10,6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8: Bullet_img = 4'd13;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//2'd2: begin
//case(angle)
//// Bullet_type_2 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd54: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd4;
//6'd26,6'd27,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd55: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd4;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd2,6'd3,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd54,6'd55,6'd56: Bullet_img = 4'd4;
//6'd53: Bullet_img = 4'd12;
//6'd4,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd15,6'd16,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd51,6'd52: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd5: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd54,6'd55,6'd56: Bullet_img = 4'd4;
//6'd53: Bullet_img = 4'd12;
//6'd4,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd15,6'd16,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd51,6'd52: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd43,6'd44,6'd55: Bullet_img = 4'd4;
//6'd52,6'd53,6'd54: Bullet_img = 4'd12;
//6'd4,6'd17,6'd24,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd18,6'd19,6'd20,6'd21,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd43,6'd44,6'd45,6'd46,6'd53,6'd54: Bullet_img = 4'd4;
//6'd52,6'd55: Bullet_img = 4'd12;
//6'd17,6'd22,6'd23: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd11,6'd14,6'd15,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd18,6'd19,6'd21,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd33,6'd34,6'd35,6'd36,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd4;
//6'd32,6'd47: Bullet_img = 4'd6;
//6'd17,6'd22,6'd23: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd7: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd21,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd32,6'd33,6'd34,6'd35,6'd36,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd4;
//6'd19,6'd31: Bullet_img = 4'd5;
//6'd18: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd7,6'd8,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd32,6'd33,6'd34,6'd35,6'd36,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd53: Bullet_img = 4'd4;
//6'd31,6'd54: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd18,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd38,6'd39,6'd40,6'd52,6'd53: Bullet_img = 4'd4;
//6'd54: Bullet_img = 4'd5;
//6'd19: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd7,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd38,6'd39,6'd40,6'd52,6'd53: Bullet_img = 4'd4;
//6'd54: Bullet_img = 4'd5;
//6'd5,6'd6,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd19: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd63,6'd64: Bullet_img = 4'd0;
//6'd53: Bullet_img = 4'd3;
//6'd20,6'd38,6'd39,6'd40,6'd52: Bullet_img = 4'd4;
//6'd54: Bullet_img = 4'd5;
//6'd4,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd19: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd2,6'd3,6'd63,6'd64: Bullet_img = 4'd0;
//6'd53: Bullet_img = 4'd3;
//6'd20,6'd52,6'd54: Bullet_img = 4'd5;
//6'd4: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd59,6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd52,6'd53: Bullet_img = 4'd3;
//6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd54: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd21,6'd22,6'd23,6'd48,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd20: Bullet_img = 4'd3;
//6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd37,6'd41,6'd42,6'd52,6'd53,6'd54: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd21,6'd22,6'd23,6'd24,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd20: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd4;
//6'd52,6'd53,6'd54: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd18,6'd21,6'd22,6'd23,6'd24,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd21,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd20,6'd55: Bullet_img = 4'd2;
//6'd54: Bullet_img = 4'd3;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd4;
//6'd52,6'd53: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd8,6'd17,6'd22,6'd23,6'd24,6'd25,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd2;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//6'd1,6'd2,6'd3,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd2;
//6'd4: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd5,6'd6,6'd13,6'd14,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd50,6'd51,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//6'd1,6'd2,6'd3,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd2;
//6'd4: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd5,6'd6,6'd14,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd50,6'd51,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd2;
//6'd4: Bullet_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd5,6'd6,6'd11,6'd12,6'd13,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//6'd1,6'd2,6'd3,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd55,6'd56: Bullet_img = 4'd2;
//6'd4: Bullet_img = 4'd13;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//6'd1,6'd2,6'd3,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd55,6'd56: Bullet_img = 4'd2;
//6'd4: Bullet_img = 4'd13;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd54: Bullet_img = 4'd14;
//6'd26,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd54: Bullet_img = 4'd4;
//6'd50: Bullet_img = 4'd8;
//6'd27,6'd28,6'd51,6'd52,6'd53: Bullet_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd8;
//6'd29,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd13;
//6'd39,6'd40: Bullet_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48: Bullet_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49: Bullet_img = 4'd4;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd4;
//6'd39,6'd40: Bullet_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd4;
//6'd47: Bullet_img = 4'd12;
//6'd37,6'd38,6'd39,6'd40,6'd45,6'd46: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44,6'd52: Bullet_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49: Bullet_img = 4'd4;
//6'd47: Bullet_img = 4'd12;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd12;
//6'd24,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd40,6'd41,6'd42,6'd43,6'd44,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd4;
//6'd47: Bullet_img = 4'd12;
//6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Bullet_img = 4'd14;
//6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd4;
//6'd47: Bullet_img = 4'd12;
//6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd4;
//6'd23,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd48,6'd49: Bullet_img = 4'd4;
//6'd50: Bullet_img = 4'd5;
//6'd43: Bullet_img = 4'd6;
//6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd50: Bullet_img = 4'd4;
//6'd51: Bullet_img = 4'd5;
//6'd21,6'd22,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd49,6'd50: Bullet_img = 4'd4;
//6'd51: Bullet_img = 4'd5;
//6'd21,6'd22,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd23,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51: Bullet_img = 4'd3;
//6'd31,6'd32,6'd40,6'd41,6'd42,6'd43,6'd49: Bullet_img = 4'd4;
//6'd52: Bullet_img = 4'd5;
//6'd20,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd44,6'd45,6'd46,6'd47,6'd48,6'd53,6'd54: Bullet_img = 4'd14;
//6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd51: Bullet_img = 4'd3;
//6'd30,6'd31,6'd32,6'd33,6'd40: Bullet_img = 4'd4;
//6'd50,6'd52: Bullet_img = 4'd5;
//6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd28,6'd29,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd60: Bullet_img = 4'd14;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51: Bullet_img = 4'd3;
//6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd52: Bullet_img = 4'd5;
//6'd24,6'd25: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53: Bullet_img = 4'd14;
//6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd37,6'd38: Bullet_img = 4'd4;
//6'd51,6'd52,6'd53: Bullet_img = 4'd5;
//6'd29: Bullet_img = 4'd6;
//6'd20,6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//6'd21,6'd22,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54: Bullet_img = 4'd14;
//6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd54: Bullet_img = 4'd2;
//6'd53: Bullet_img = 4'd3;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd51,6'd52: Bullet_img = 4'd5;
//6'd21,6'd23: Bullet_img = 4'd13;
//6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd53,6'd54,6'd55: Bullet_img = 4'd2;
//6'd30,6'd31,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd29,6'd51,6'd52: Bullet_img = 4'd5;
//6'd13: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd32,6'd33,6'd34,6'd35,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd14,6'd15,6'd16,6'd17,6'd18,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd2;
//6'd8,6'd9,6'd10,6'd12,6'd13,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd56,6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd15,6'd16,6'd17,6'd18,6'd19,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd40,6'd41: Bullet_img = 4'd5;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd12,6'd13,6'd14,6'd20,6'd21: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd16,6'd17,6'd19,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd54,6'd55,6'd56,6'd57: Bullet_img = 4'd2;
//6'd18,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd4;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd15: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd14,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd16,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd56,6'd57: Bullet_img = 4'd2;
//6'd18,6'd19,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd4;
//6'd17,6'd37: Bullet_img = 4'd5;
//6'd2,6'd3,6'd5,6'd6,6'd7,6'd8,6'd15: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd12,6'd13,6'd43,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd2,6'd6: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd9,6'd17,6'd41,6'd42,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd55,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19,6'd37: Bullet_img = 4'd4;
//6'd2,6'd18: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd4,6'd54,6'd55,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd57: Bullet_img = 4'd4;
//6'd2,6'd19: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd37,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd52,6'd53,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd5;
//6'd19,6'd54,6'd55,6'd56: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd6,6'd7,6'd23,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd7,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd3;
//6'd53: Bullet_img = 4'd8;
//6'd13: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd6,6'd22,6'd23,6'd24,6'd25,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd3;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd13;
//6'd8,6'd9,6'd14,6'd15,6'd16,6'd17,6'd20,6'd27,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd21: Bullet_img = 4'd2;
//6'd8,6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd35,6'd36: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd23,6'd24,6'd25,6'd26,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd1;
//6'd22: Bullet_img = 4'd2;
//6'd6,6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd13;
//6'd11,6'd12,6'd18,6'd19: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd16,6'd17,6'd18: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd19,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd5: Bullet_img = 4'd13;
//6'd6,6'd7,6'd10,6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd14;
//6'd18,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd14;
//6'd17,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36: Bullet_img = 4'd8;
//6'd32,6'd33: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd14;
//6'd11,6'd16,6'd17,6'd30,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd4;
//6'd32: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd14;
//6'd9,6'd10,6'd11,6'd17,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd14;
//6'd9,6'd10,6'd15,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd14;
//6'd9,6'd10: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8: Bullet_img = 4'd13;
//6'd11: Bullet_img = 4'd14;
//6'd9,6'd10,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9: Bullet_img = 4'd13;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45,6'd46: Bullet_img = 4'd13;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46,6'd47: Bullet_img = 4'd13;
//6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48: Bullet_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd42,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd42,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd53: Bullet_img = 4'd13;
//6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd41,6'd42,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd53: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52: Bullet_img = 4'd14;
//6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd53: Bullet_img = 4'd13;
//6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52: Bullet_img = 4'd14;
//6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd51,6'd52,6'd53: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd49,6'd50: Bullet_img = 4'd14;
//6'd41,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd49: Bullet_img = 4'd14;
//6'd41,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd48,6'd52: Bullet_img = 4'd14;
//6'd40,6'd41,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd58,6'd59: Bullet_img = 4'd13;
//6'd41,6'd42,6'd43,6'd47,6'd51,6'd52,6'd53,6'd55,6'd56: Bullet_img = 4'd14;
//6'd44,6'd45,6'd46,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28: Bullet_img = 4'd4;
//6'd27,6'd47,6'd48,6'd49,6'd59,6'd60: Bullet_img = 4'd13;
//6'd41,6'd42,6'd46,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd14;
//6'd43,6'd44,6'd45,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39: Bullet_img = 4'd1;
//6'd26,6'd27,6'd47,6'd48: Bullet_img = 4'd13;
//6'd45,6'd46,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd14;
//6'd25,6'd40,6'd41,6'd42,6'd43,6'd44,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd1;
//6'd38,6'd39: Bullet_img = 4'd2;
//6'd56,6'd59: Bullet_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd57,6'd58: Bullet_img = 4'd14;
//6'd28,6'd29,6'd30,6'd32,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39: Bullet_img = 4'd2;
//6'd40: Bullet_img = 4'd3;
//6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd13;
//6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54: Bullet_img = 4'd14;
//6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd38,6'd42,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41: Bullet_img = 4'd3;
//6'd54,6'd55,6'd56,6'd57: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42: Bullet_img = 4'd4;
//6'd41: Bullet_img = 4'd5;
//6'd43,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd13;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51,6'd52: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd4;
//6'd44,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd13;
//6'd34,6'd35,6'd36,6'd40,6'd41,6'd47,6'd48,6'd51: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd37,6'd38,6'd39,6'd45,6'd46,6'd49,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44: Bullet_img = 4'd4;
//6'd46,6'd48,6'd51,6'd53,6'd54: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd45,6'd50,6'd52: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45: Bullet_img = 4'd4;
//6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd4;
//6'd44: Bullet_img = 4'd12;
//6'd51: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44,6'd45: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27: Bullet_img = 4'd4;
//6'd44: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd4;
//6'd45: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd28,6'd36: Bullet_img = 4'd5;
//6'd42: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd35,6'd36: Bullet_img = 4'd4;
//6'd37: Bullet_img = 4'd5;
//6'd41,6'd42,6'd46: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd40,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd10,6'd13,6'd14,6'd15,6'd16,6'd17,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd47: Bullet_img = 4'd4;
//6'd37: Bullet_img = 4'd6;
//6'd11: Bullet_img = 4'd8;
//6'd10,6'd41,6'd42,6'd43,6'd46: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd39,6'd40,6'd44,6'd45: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd29,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd4;
//6'd25: Bullet_img = 4'd5;
//6'd9,6'd10,6'd40,6'd41,6'd42,6'd46: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd28,6'd30,6'd31,6'd32,6'd38,6'd39,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd4;
//6'd24: Bullet_img = 4'd5;
//6'd9,6'd39,6'd40,6'd41,6'd42,6'd46: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd31,6'd32,6'd38,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd4;
//6'd40,6'd41: Bullet_img = 4'd13;
//6'd9,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd35,6'd36: Bullet_img = 4'd4;
//6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd12,6'd14: Bullet_img = 4'd2;
//6'd39,6'd40,6'd41: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd10,6'd11,6'd13,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd2;
//6'd38,6'd39,6'd40,6'd45,6'd46: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd2;
//6'd27,6'd28: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd5;
//6'd38,6'd39,6'd40,6'd41,6'd45,6'd46: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14: Bullet_img = 4'd2;
//6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd4;
//6'd15,6'd16,6'd17: Bullet_img = 4'd5;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd2;
//6'd14,6'd18: Bullet_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd15,6'd16,6'd17: Bullet_img = 4'd5;
//6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33,6'd34,6'd35,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd3;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd15,6'd16,6'd18,6'd19: Bullet_img = 4'd5;
//6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd13;
//6'd14,6'd20,6'd21,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd3;
//6'd19,6'd20,6'd28: Bullet_img = 4'd4;
//6'd16,6'd17: Bullet_img = 4'd5;
//6'd26: Bullet_img = 4'd6;
//6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd13;
//6'd15,6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd4;
//6'd17,6'd18: Bullet_img = 4'd5;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd13;
//6'd15,6'd16,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22: Bullet_img = 4'd4;
//6'd18,6'd19: Bullet_img = 4'd5;
//6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd19,6'd20: Bullet_img = 4'd5;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//6'd9,6'd14,6'd15,6'd16,6'd17,6'd18,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd5;
//6'd23,6'd24: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd25,6'd26,6'd27,6'd28,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd24: Bullet_img = 4'd12;
//6'd25,6'd26,6'd28,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd27,6'd29,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd4;
//6'd21,6'd23,6'd24: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27,6'd32: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24: Bullet_img = 4'd4;
//6'd25: Bullet_img = 4'd12;
//6'd26: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd4;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34: Bullet_img = 4'd14;
//6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd4;
//6'd15,6'd16,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd14;
//6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27: Bullet_img = 4'd13;
//6'd25,6'd26,6'd28: Bullet_img = 4'd14;
//6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27: Bullet_img = 4'd13;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35: Bullet_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37: Bullet_img = 4'd13;
//6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44: Bullet_img = 4'd13;
//6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd32,6'd33,6'd34,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd43,6'd44: Bullet_img = 4'd14;
//6'd32,6'd33,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd13;
//6'd34,6'd35,6'd36,6'd39,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd32,6'd33,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd51,6'd52: Bullet_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44,6'd53: Bullet_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd42,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//6'd33,6'd39,6'd40,6'd41,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43,6'd53: Bullet_img = 4'd13;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd44,6'd45,6'd46,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//6'd33,6'd39,6'd40,6'd47,6'd48,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43,6'd53: Bullet_img = 4'd13;
//6'd35,6'd36,6'd37,6'd38,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd33,6'd34,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd35,6'd36,6'd37,6'd40,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd34,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd36,6'd37,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd35,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd35,6'd36,6'd40,6'd43,6'd44,6'd45,6'd46,6'd48: Bullet_img = 4'd14;
//6'd34,6'd37,6'd38,6'd39,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd35,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34: Bullet_img = 4'd1;
//6'd48,6'd49,6'd50: Bullet_img = 4'd13;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47: Bullet_img = 4'd14;
//6'd35,6'd36,6'd37,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd1;
//6'd34: Bullet_img = 4'd2;
//6'd50: Bullet_img = 4'd13;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd3;
//6'd37: Bullet_img = 4'd5;
//6'd39,6'd44,6'd47,6'd48: Bullet_img = 4'd13;
//6'd38,6'd40,6'd41,6'd43,6'd46: Bullet_img = 4'd14;
//6'd34,6'd42,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd38,6'd39: Bullet_img = 4'd4;
//6'd37,6'd42: Bullet_img = 4'd5;
//6'd40,6'd43,6'd45,6'd46,6'd48: Bullet_img = 4'd13;
//6'd41: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41: Bullet_img = 4'd4;
//6'd42: Bullet_img = 4'd5;
//6'd23: Bullet_img = 4'd13;
//6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd24,6'd26,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd4;
//6'd22: Bullet_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd21,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd8;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47: Bullet_img = 4'd4;
//6'd42,6'd46: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd47: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37: Bullet_img = 4'd5;
//6'd41,6'd42,6'd43,6'd47: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37: Bullet_img = 4'd4;
//6'd38: Bullet_img = 4'd5;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd36,6'd37: Bullet_img = 4'd4;
//6'd38: Bullet_img = 4'd6;
//6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd41,6'd42,6'd43,6'd44,6'd48: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd40,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd29: Bullet_img = 4'd5;
//6'd42,6'd43,6'd44,6'd48,6'd49: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd42,6'd43,6'd44,6'd48,6'd49: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd31,6'd32,6'd33,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd30,6'd34,6'd35,6'd36,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd28,6'd29,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd27: Bullet_img = 4'd5;
//6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd27: Bullet_img = 4'd5;
//6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd4;
//6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd8;
//6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd13,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd8;
//6'd13,6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd13,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd4;
//6'd13,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd13,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd35,6'd36,6'd37,6'd38,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd32: Bullet_img = 4'd6;
//6'd39,6'd40,6'd41: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd15,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd21,6'd22,6'd23: Bullet_img = 4'd5;
//6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd24: Bullet_img = 4'd3;
//6'd21,6'd22,6'd23,6'd25: Bullet_img = 4'd5;
//6'd38,6'd39,6'd40: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd18,6'd19,6'd20: Bullet_img = 4'd2;
//6'd24,6'd25: Bullet_img = 4'd3;
//6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd21,6'd22,6'd23: Bullet_img = 4'd5;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd23,6'd24,6'd25: Bullet_img = 4'd5;
//6'd36: Bullet_img = 4'd13;
//6'd21,6'd22,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd26,6'd27: Bullet_img = 4'd5;
//6'd31,6'd32,6'd33: Bullet_img = 4'd12;
//6'd34,6'd35,6'd36: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd28: Bullet_img = 4'd5;
//6'd32: Bullet_img = 4'd12;
//6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd35: Bullet_img = 4'd4;
//6'd32,6'd33,6'd34: Bullet_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd4;
//6'd30: Bullet_img = 4'd12;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd37: Bullet_img = 4'd13;
//6'd18,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd36: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34: Bullet_img = 4'd4;
//6'd36: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd35: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd33,6'd34,6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd44: Bullet_img = 4'd13;
//6'd33,6'd34,6'd41,6'd42: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd44: Bullet_img = 4'd13;
//6'd33,6'd34,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd44: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd33,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd23,6'd24,6'd28,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd36,6'd37,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd23,6'd24,6'd28,6'd29,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd23,6'd24,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd23,6'd24,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd36,6'd37,6'd38,6'd39,6'd41: Bullet_img = 4'd14;
//6'd25,6'd31,6'd32,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd25,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd26,6'd28,6'd29,6'd30,6'd33,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd25,6'd27,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd26,6'd27,6'd31,6'd32,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41: Bullet_img = 4'd14;
//6'd28,6'd31,6'd32,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd29,6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd41: Bullet_img = 4'd14;
//6'd28,6'd31,6'd32,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40,6'd41: Bullet_img = 4'd13;
//6'd30,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd29,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31: Bullet_img = 4'd1;
//6'd38: Bullet_img = 4'd5;
//6'd34,6'd35,6'd36: Bullet_img = 4'd13;
//6'd32,6'd33,6'd37: Bullet_img = 4'd14;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd2;
//6'd31,6'd32: Bullet_img = 4'd3;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd33: Bullet_img = 4'd5;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd4;
//6'd45: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd4;
//6'd41,6'd46: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd41,6'd46,6'd47: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd48: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43,6'd44,6'd49,6'd50: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd5;
//6'd19: Bullet_img = 4'd8;
//6'd42,6'd43,6'd44,6'd45,6'd49,6'd50: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd4;
//6'd39: Bullet_img = 4'd6;
//6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd44,6'd45: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd4;
//6'd31: Bullet_img = 4'd5;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd4;
//6'd31: Bullet_img = 4'd5;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd4;
//6'd31: Bullet_img = 4'd5;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd4;
//6'd39: Bullet_img = 4'd6;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd8;
//6'd44: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28: Bullet_img = 4'd2;
//6'd32: Bullet_img = 4'd3;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd29,6'd30,6'd31,6'd33: Bullet_img = 4'd5;
//6'd40,6'd41: Bullet_img = 4'd12;
//6'd20,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd2;
//6'd32,6'd33,6'd34: Bullet_img = 4'd3;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd44: Bullet_img = 4'd4;
//6'd29,6'd30,6'd31: Bullet_img = 4'd5;
//6'd41,6'd42,6'd43: Bullet_img = 4'd12;
//6'd20: Bullet_img = 4'd13;
//6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd2;
//6'd29: Bullet_img = 4'd3;
//6'd20,6'd38,6'd39,6'd40,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd5;
//6'd41: Bullet_img = 4'd12;
//6'd47: Bullet_img = 4'd13;
//6'd21,6'd45,6'd46: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd2;
//6'd38,6'd39,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd40: Bullet_img = 4'd12;
//6'd46: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd45: Bullet_img = 4'd14;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25: Bullet_img = 4'd2;
//6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd37,6'd38: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd13;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd13;
//6'd29,6'd30: Bullet_img = 4'd14;
//6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd32,6'd33: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd13;
//6'd22,6'd23,6'd29,6'd30: Bullet_img = 4'd14;
//6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd32,6'd33,6'd34: Bullet_img = 4'd13;
//6'd22,6'd23,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd24,6'd25,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd24,6'd25,6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd32: Bullet_img = 4'd14;
//6'd15,6'd16,6'd17,6'd18,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd20,6'd21,6'd24,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd13,6'd14,6'd18,6'd19,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd34,6'd35: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd24,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd22,6'd23,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd34,6'd35,6'd36: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd25,6'd28,6'd29,6'd30,6'd31,6'd33: Bullet_img = 4'd14;
//6'd14,6'd15,6'd22,6'd23,6'd24,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd14,6'd15,6'd23,6'd24,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//6'd15,6'd17,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd20,6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//6'd17,6'd19,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd5;
//6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd24,6'd25,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33: Bullet_img = 4'd4;
//6'd30: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd31: Bullet_img = 4'd14;
//6'd21,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32: Bullet_img = 4'd4;
//6'd28,6'd29,6'd35: Bullet_img = 4'd13;
//6'd24,6'd27: Bullet_img = 4'd14;
//6'd23,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd1;
//6'd27: Bullet_img = 4'd3;
//6'd29,6'd42: Bullet_img = 4'd4;
//6'd28: Bullet_img = 4'd5;
//6'd34,6'd35,6'd38,6'd41: Bullet_img = 4'd13;
//6'd26,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd1;
//6'd25: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd3;
//6'd34,6'd35,6'd37,6'd42,6'd43: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd2;
//6'd42,6'd43: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40,6'd47,6'd48: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37: Bullet_img = 4'd4;
//6'd36: Bullet_img = 4'd5;
//6'd38: Bullet_img = 4'd6;
//6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd41,6'd42,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd19,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd18,6'd19,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd42,6'd43,6'd44,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd19,6'd46,6'd47,6'd48: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44,6'd45,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd18,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd8;
//6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd33,6'd34,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd32: Bullet_img = 4'd5;
//6'd48,6'd49,6'd50: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd44: Bullet_img = 4'd4;
//6'd48,6'd49,6'd50: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd34,6'd36,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd35,6'd36,6'd37,6'd38,6'd39,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd49: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd49: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd41,6'd42,6'd43: Bullet_img = 4'd4;
//6'd44: Bullet_img = 4'd6;
//6'd49: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42: Bullet_img = 4'd4;
//6'd49: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd54: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd51: Bullet_img = 4'd4;
//6'd46,6'd47,6'd49,6'd50: Bullet_img = 4'd12;
//6'd48: Bullet_img = 4'd13;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd52,6'd53: Bullet_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51: Bullet_img = 4'd4;
//6'd48: Bullet_img = 4'd12;
//6'd53: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd52: Bullet_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd4;
//6'd48: Bullet_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd41: Bullet_img = 4'd3;
//6'd42,6'd43,6'd45,6'd46,6'd47,6'd50,6'd51: Bullet_img = 4'd4;
//6'd40,6'd44: Bullet_img = 4'd5;
//6'd48: Bullet_img = 4'd12;
//6'd32,6'd35,6'd36,6'd37,6'd38,6'd49: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40,6'd41: Bullet_img = 4'd3;
//6'd46: Bullet_img = 4'd4;
//6'd36,6'd37,6'd38,6'd42,6'd43: Bullet_img = 4'd5;
//6'd35,6'd44,6'd45,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35: Bullet_img = 4'd2;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd5;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd37: Bullet_img = 4'd3;
//6'd38: Bullet_img = 4'd5;
//6'd27: Bullet_img = 4'd8;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd26,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd2;
//6'd28: Bullet_img = 4'd13;
//6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd2;
//6'd28: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd31,6'd32,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd28: Bullet_img = 4'd13;
//6'd29,6'd30,6'd42,6'd47,6'd48: Bullet_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34: Bullet_img = 4'd2;
//6'd29: Bullet_img = 4'd4;
//6'd47: Bullet_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd14;
//6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd21: Bullet_img = 4'd13;
//6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd22: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21: Bullet_img = 4'd14;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21: Bullet_img = 4'd14;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20: Bullet_img = 4'd14;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd14;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd18,6'd20,6'd21,6'd23: Bullet_img = 4'd14;
//6'd19,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd15,6'd25,6'd27: Bullet_img = 4'd13;
//6'd13,6'd14,6'd17,6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd26: Bullet_img = 4'd14;
//6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//6'd13,6'd14,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd18,6'd27: Bullet_img = 4'd13;
//6'd14,6'd15,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26: Bullet_img = 4'd14;
//6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd27: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd14;
//6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7,6'd8,6'd18,6'd19,6'd20,6'd26: Bullet_img = 4'd13;
//6'd13,6'd14,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd14;
//6'd10,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36: Bullet_img = 4'd4;
//6'd6,6'd7,6'd19,6'd20: Bullet_img = 4'd13;
//6'd13,6'd14,6'd17,6'd18,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd14;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd15,6'd16: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd5,6'd6,6'd26,6'd35,6'd36,6'd37,6'd38,6'd42,6'd43: Bullet_img = 4'd13;
//6'd10,6'd13,6'd14,6'd15,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd39: Bullet_img = 4'd14;
//6'd7,6'd8,6'd9,6'd11,6'd12,6'd16,6'd17,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd4;
//6'd5,6'd30,6'd33,6'd42,6'd43: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44: Bullet_img = 4'd14;
//6'd6,6'd7,6'd8,6'd17,6'd18,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd4;
//6'd28: Bullet_img = 4'd12;
//6'd25,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd6,6'd7,6'd8,6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd4;
//6'd24,6'd30,6'd36: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd7,6'd8,6'd9,6'd19,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25: Bullet_img = 4'd4;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Bullet_img = 4'd13;
//6'd13,6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd14,6'd20,6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd5;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd43,6'd44: Bullet_img = 4'd13;
//6'd14,6'd18,6'd19,6'd22,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd42,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd9,6'd12,6'd13,6'd15,6'd16,6'd17,6'd20,6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd1;
//6'd22,6'd23: Bullet_img = 4'd3;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd13,6'd17,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd1;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd2;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd35: Bullet_img = 4'd5;
//6'd36: Bullet_img = 4'd6;
//6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42,6'd43,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd41,6'd42,6'd43,6'd44,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd4;
//6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd54: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd45,6'd46: Bullet_img = 4'd4;
//6'd51,6'd52: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd44,6'd45,6'd46: Bullet_img = 4'd4;
//6'd51: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd47,6'd48,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd36,6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd52: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd35,6'd37,6'd40,6'd41,6'd42,6'd48,6'd49,6'd50,6'd51,6'd53,6'd54,6'd55,6'd56,6'd57: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd4;
//6'd19,6'd20,6'd53,6'd57,6'd58: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd38,6'd39,6'd40,6'd41,6'd42,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd44,6'd45,6'd46: Bullet_img = 4'd4;
//6'd47: Bullet_img = 4'd6;
//6'd20,6'd52,6'd53,6'd54: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd48,6'd49,6'd50,6'd51,6'd55,6'd56,6'd57: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd45,6'd46,6'd55: Bullet_img = 4'd4;
//6'd37: Bullet_img = 4'd5;
//6'd54: Bullet_img = 4'd12;
//6'd52,6'd53: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd56,6'd57: Bullet_img = 4'd14;
//6'd20,6'd23,6'd24,6'd25,6'd26,6'd27,6'd32,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37,6'd54,6'd55,6'd56: Bullet_img = 4'd4;
//6'd38: Bullet_img = 4'd5;
//6'd51,6'd52,6'd53: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31,6'd32,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd50,6'd52,6'd54,6'd55,6'd56: Bullet_img = 4'd4;
//6'd51,6'd53: Bullet_img = 4'd12;
//6'd30,6'd31,6'd32,6'd33,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd4;
//6'd31,6'd32,6'd33,6'd34,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd4;
//6'd53: Bullet_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47,6'd54,6'd55: Bullet_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd36,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48,6'd49,6'd52: Bullet_img = 4'd4;
//6'd50,6'd51: Bullet_img = 4'd5;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48: Bullet_img = 4'd4;
//6'd46,6'd49,6'd50: Bullet_img = 4'd5;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45,6'd46,6'd47: Bullet_img = 4'd3;
//6'd48,6'd49: Bullet_img = 4'd5;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd3;
//6'd44,6'd45,6'd47,6'd48: Bullet_img = 4'd5;
//6'd36,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd5;
//6'd39,6'd40,6'd41,6'd42,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd2;
//6'd44,6'd45,6'd46: Bullet_img = 4'd5;
//6'd47,6'd48,6'd50,6'd51,6'd55,6'd56: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd49,6'd52,6'd53,6'd54,6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd2;
//6'd45: Bullet_img = 4'd3;
//6'd46: Bullet_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd2;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd2;
//6'd33,6'd37,6'd38,6'd39,6'd40,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd2;
//6'd36: Bullet_img = 4'd8;
//6'd38,6'd39,6'd40,6'd41,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd2;
//6'd36,6'd37: Bullet_img = 4'd13;
//6'd35,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42: Bullet_img = 4'd2;
//6'd37,6'd38: Bullet_img = 4'd13;
//6'd39,6'd50: Bullet_img = 4'd14;
//6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd4;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12: Bullet_img = 4'd13;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd13,6'd14,6'd15: Bullet_img = 4'd13;
//6'd12: Bullet_img = 4'd14;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12: Bullet_img = 4'd14;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18,6'd20,6'd37: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd19: Bullet_img = 4'd14;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd20,6'd21,6'd35,6'd36,6'd37: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd18,6'd19,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd11: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30: Bullet_img = 4'd4;
//6'd20,6'd21,6'd31,6'd32: Bullet_img = 4'd13;
//6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd11,6'd12,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd20,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7,6'd8,6'd21,6'd39: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd6,6'd7,6'd9,6'd11,6'd20,6'd28,6'd35,6'd36,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd8,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd37,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//endcase
//end
//6'd20: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd22,6'd24,6'd25,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd4;
//6'd10,6'd11,6'd12,6'd13,6'd21,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//endcase
//end
//6'd21: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd24,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd23: Bullet_img = 4'd4;
//6'd22: Bullet_img = 4'd5;
//default: Bullet_img = 4'd13;
//6'd9,6'd10,6'd16,6'd17,6'd18,6'd19,6'd27,6'd28,6'd29,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd20,6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd4;
//6'd14,6'd15,6'd32,6'd34,6'd35,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd4;
//6'd21,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd21,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd20,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd21,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd6;
//6'd4,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8,6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd21: Bullet_img = 4'd5;
//6'd3,6'd50,6'd51: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd4,6'd5,6'd6,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd20: Bullet_img = 4'd3;
//6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd4;
//6'd3,6'd51,6'd52,6'd53,6'd58: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd4,6'd5,6'd18,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd1;
//6'd20: Bullet_img = 4'd3;
//6'd36,6'd37,6'd45,6'd46,6'd55: Bullet_img = 4'd4;
//6'd3,6'd53,6'd54: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd4,6'd5,6'd17,6'd18,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd17,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd1;
//6'd19: Bullet_img = 4'd2;
//6'd44,6'd45,6'd46,6'd47,6'd55,6'd56,6'd57: Bullet_img = 4'd4;
//6'd53,6'd54: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6,6'd12,6'd13,6'd14,6'd15,6'd16,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd38,6'd39,6'd44,6'd45,6'd46,6'd47,6'd56,6'd57,6'd58: Bullet_img = 4'd4;
//6'd54,6'd55: Bullet_img = 4'd12;
//6'd53: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40,6'd44,6'd45,6'd46,6'd47,6'd56,6'd57: Bullet_img = 4'd4;
//6'd48: Bullet_img = 4'd6;
//6'd53,6'd54,6'd55: Bullet_img = 4'd12;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd7,6'd8,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40,6'd45,6'd46,6'd47,6'd53,6'd54,6'd56: Bullet_img = 4'd4;
//6'd55: Bullet_img = 4'd12;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd51,6'd52,6'd57: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd4;
//default: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd4;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36,6'd37,6'd38,6'd51,6'd52,6'd53: Bullet_img = 4'd4;
//6'd39,6'd54: Bullet_img = 4'd5;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd51,6'd52: Bullet_img = 4'd4;
//6'd40,6'd53: Bullet_img = 4'd5;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd50,6'd51,6'd52: Bullet_img = 4'd4;
//6'd53: Bullet_img = 4'd5;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd41,6'd42,6'd43,6'd44,6'd45,6'd47,6'd48,6'd49,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd46,6'd61: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd51: Bullet_img = 4'd3;
//6'd39,6'd40: Bullet_img = 4'd4;
//6'd50,6'd52: Bullet_img = 4'd5;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd36,6'd37,6'd38,6'd60,6'd61: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51: Bullet_img = 4'd3;
//6'd52: Bullet_img = 4'd5;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd39,6'd40,6'd57,6'd58,6'd59,6'd60,6'd61: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd4;
//6'd49,6'd50,6'd51: Bullet_img = 4'd5;
//6'd22: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51: Bullet_img = 4'd5;
//6'd23: Bullet_img = 4'd13;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd52,6'd53: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd5;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd2;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd2;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd2;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50: Bullet_img = 4'd2;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51: Bullet_img = 4'd2;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50: Bullet_img = 4'd2;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd13;
//6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45,6'd46: Bullet_img = 4'd13;
//6'd47: Bullet_img = 4'd14;
//6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37: Bullet_img = 4'd13;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37: Bullet_img = 4'd13;
//6'd36,6'd38,6'd39: Bullet_img = 4'd14;
//6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41: Bullet_img = 4'd4;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd44,6'd45,6'd46,6'd48,6'd49: Bullet_img = 4'd14;
//6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd4;
//6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41,6'd42: Bullet_img = 4'd4;
//6'd39: Bullet_img = 4'd12;
//6'd38: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42: Bullet_img = 4'd4;
//6'd40,6'd41,6'd43: Bullet_img = 4'd12;
//6'd32,6'd37,6'd38,6'd39: Bullet_img = 4'd13;
//6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd40: Bullet_img = 4'd12;
//6'd31,6'd32,6'd33,6'd34,6'd36,6'd38,6'd39: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd35,6'd37,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43: Bullet_img = 4'd4;
//6'd44: Bullet_img = 4'd5;
//6'd40,6'd41: Bullet_img = 4'd12;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd36,6'd37,6'd38,6'd39,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42,6'd43: Bullet_img = 4'd4;
//6'd44,6'd45: Bullet_img = 4'd5;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd46,6'd47,6'd48,6'd49,6'd55: Bullet_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd43,6'd44: Bullet_img = 4'd4;
//6'd45,6'd46: Bullet_img = 4'd5;
//6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd47,6'd48: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd44,6'd45: Bullet_img = 4'd4;
//6'd46,6'd47: Bullet_img = 4'd5;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd48,6'd49: Bullet_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd3;
//6'd36,6'd44,6'd45: Bullet_img = 4'd4;
//6'd47,6'd48: Bullet_img = 4'd5;
//6'd38: Bullet_img = 4'd6;
//6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd31,6'd32,6'd33,6'd34,6'd35,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43,6'd49: Bullet_img = 4'd14;
//6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46,6'd47: Bullet_img = 4'd3;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd45,6'd48,6'd49: Bullet_img = 4'd5;
//6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd40,6'd41,6'd42,6'd43,6'd44,6'd50: Bullet_img = 4'd14;
//6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd51: Bullet_img = 4'd2;
//6'd46,6'd50: Bullet_img = 4'd3;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd47,6'd48,6'd49: Bullet_img = 4'd5;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51,6'd52: Bullet_img = 4'd2;
//6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd47,6'd48,6'd49: Bullet_img = 4'd5;
//6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd2;
//6'd36,6'd37: Bullet_img = 4'd4;
//6'd48: Bullet_img = 4'd5;
//6'd18,6'd19,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd2;
//6'd18,6'd19,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd52,6'd55: Bullet_img = 4'd2;
//6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd49,6'd51,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd35: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd56: Bullet_img = 4'd4;
//6'd23,6'd24: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd25,6'd26,6'd31,6'd32,6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd55: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd36,6'd56: Bullet_img = 4'd4;
//6'd40: Bullet_img = 4'd5;
//6'd18,6'd22,6'd23,6'd24,6'd25,6'd55: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd26,6'd32,6'd33,6'd37,6'd38,6'd39,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd35,6'd37,6'd38,6'd40,6'd41,6'd42: Bullet_img = 4'd4;
//6'd39: Bullet_img = 4'd5;
//6'd18,6'd22,6'd23,6'd24,6'd54,6'd55: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd32,6'd33,6'd34,6'd36,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd4;
//6'd27: Bullet_img = 4'd6;
//6'd53: Bullet_img = 4'd8;
//6'd18,6'd21,6'd22,6'd23,6'd54: Bullet_img = 4'd13;
//6'd19,6'd20,6'd24,6'd25,6'd26,6'd31,6'd32,6'd33,6'd34,6'd35,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd14;
//6'd42,6'd43,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd4;
//6'd27: Bullet_img = 4'd5;
//6'd18,6'd22,6'd23: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd24,6'd25,6'd26,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd41,6'd42,6'd47,6'd48,6'd49,6'd50,6'd51,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39: Bullet_img = 4'd4;
//6'd28,6'd36: Bullet_img = 4'd5;
//6'd22: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd40,6'd41,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd4;
//6'd19: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd39,6'd40,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd38,6'd39,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd38,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd12;
//6'd13: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd4;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd4;
//6'd10,6'd11,6'd13,6'd16,6'd18: Bullet_img = 4'd13;
//6'd12,6'd14,6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//6'd15,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd4;
//6'd9,6'd10,6'd11,6'd12,6'd20: Bullet_img = 4'd13;
//6'd13,6'd16,6'd17,6'd23,6'd24,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd14,6'd15,6'd18,6'd19,6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd4;
//6'd23: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd11,6'd21: Bullet_img = 4'd13;
//6'd12,6'd13,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd14;
//6'd14,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd3;
//6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd2;
//6'd24: Bullet_img = 4'd3;
//6'd6,6'd7,6'd8,6'd9: Bullet_img = 4'd13;
//6'd10,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd23: Bullet_img = 4'd14;
//6'd11,6'd12,6'd22,6'd26,6'd27,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd1;
//6'd25,6'd26: Bullet_img = 4'd2;
//6'd5,6'd8: Bullet_img = 4'd13;
//6'd6,6'd7,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd14;
//6'd21,6'd22,6'd23,6'd32,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25: Bullet_img = 4'd1;
//6'd16,6'd17,6'd37,6'd38: Bullet_img = 4'd13;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd18,6'd19: Bullet_img = 4'd14;
//6'd5,6'd20,6'd21,6'd22,6'd23,6'd24,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36: Bullet_img = 4'd4;
//6'd4,6'd5,6'd15,6'd16,6'd17,6'd37: Bullet_img = 4'd13;
//6'd6,6'd7,6'd8,6'd9,6'd10,6'd12,6'd13,6'd14,6'd18,6'd22,6'd23: Bullet_img = 4'd14;
//6'd11,6'd19,6'd20,6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd5,6'd6,6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd8,6'd9,6'd11,6'd12,6'd13,6'd17,6'd21,6'd22,6'd23: Bullet_img = 4'd14;
//6'd10,6'd18,6'd19,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15: Bullet_img = 4'd13;
//6'd12,6'd16,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14: Bullet_img = 4'd13;
//6'd15,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd16,6'd17,6'd18,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13: Bullet_img = 4'd13;
//6'd14,6'd15,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd16,6'd17,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd13;
//6'd12,6'd13,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd23: Bullet_img = 4'd14;
//6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd13;
//6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd23,6'd24: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21: Bullet_img = 4'd14;
//6'd17,6'd18,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21: Bullet_img = 4'd14;
//6'd17,6'd18,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd14;
//6'd16,6'd17,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd14;
//6'd17,6'd18,6'd21,6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18: Bullet_img = 4'd13;
//6'd19,6'd20: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19: Bullet_img = 4'd13;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31: Bullet_img = 4'd4;
//6'd28: Bullet_img = 4'd13;
//6'd29,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32: Bullet_img = 4'd4;
//6'd27: Bullet_img = 4'd13;
//6'd28,6'd29,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd46: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd30,6'd31,6'd32: Bullet_img = 4'd12;
//6'd26,6'd27,6'd28,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35: Bullet_img = 4'd4;
//6'd36: Bullet_img = 4'd5;
//6'd32: Bullet_img = 4'd12;
//6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd37,6'd38: Bullet_img = 4'd5;
//6'd31,6'd32,6'd33: Bullet_img = 4'd12;
//6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd39,6'd40,6'd41: Bullet_img = 4'd5;
//6'd28: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd42,6'd43: Bullet_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45,6'd46,6'd48: Bullet_img = 4'd2;
//6'd39,6'd40: Bullet_img = 4'd3;
//6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd41,6'd42,6'd43: Bullet_img = 4'd5;
//6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd2;
//6'd40: Bullet_img = 4'd3;
//6'd39,6'd41,6'd42,6'd43: Bullet_img = 4'd5;
//6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47,6'd49: Bullet_img = 4'd2;
//6'd41,6'd42,6'd43: Bullet_img = 4'd5;
//6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd2;
//6'd32: Bullet_img = 4'd6;
//6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd52: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd51: Bullet_img = 4'd14;
//6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24,6'd51: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd28,6'd34,6'd35,6'd36,6'd37,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd38,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd22,6'd23,6'd24,6'd51: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32: Bullet_img = 4'd4;
//6'd50: Bullet_img = 4'd8;
//6'd21,6'd22,6'd23,6'd51: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd4;
//6'd50: Bullet_img = 4'd8;
//6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39: Bullet_img = 4'd4;
//6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd38,6'd39: Bullet_img = 4'd4;
//6'd37: Bullet_img = 4'd5;
//6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd40,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd33,6'd35,6'd36,6'd38,6'd39: Bullet_img = 4'd4;
//6'd37: Bullet_img = 4'd5;
//6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd40,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd31,6'd32,6'd33,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd21,6'd22: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd23,6'd24,6'd28,6'd29,6'd30,6'd34,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd39,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd4;
//6'd15,6'd16,6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd36,6'd37: Bullet_img = 4'd4;
//6'd35: Bullet_img = 4'd5;
//6'd15,6'd16,6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd38,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd36,6'd37: Bullet_img = 4'd4;
//6'd16,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd38,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd37: Bullet_img = 4'd4;
//6'd26: Bullet_img = 4'd6;
//6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd38,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd4;
//6'd26: Bullet_img = 4'd5;
//6'd21,6'd22: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd23,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27: Bullet_img = 4'd5;
//6'd17,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd24,6'd25,6'd26,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd22: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd4;
//6'd18,6'd22: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd8;
//6'd21,6'd22: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd31: Bullet_img = 4'd14;
//6'd30,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd4;
//6'd42: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24: Bullet_img = 4'd4;
//6'd22: Bullet_img = 4'd5;
//6'd41: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27: Bullet_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36,6'd38,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd41: Bullet_img = 4'd4;
//6'd22,6'd27: Bullet_img = 4'd5;
//6'd16,6'd18,6'd19,6'd21,6'd24: Bullet_img = 4'd13;
//6'd23: Bullet_img = 4'd14;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd3;
//6'd27: Bullet_img = 4'd5;
//6'd16,6'd17,6'd20,6'd25: Bullet_img = 4'd13;
//6'd18,6'd21,6'd23,6'd24,6'd26: Bullet_img = 4'd14;
//6'd19,6'd22,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29: Bullet_img = 4'd1;
//6'd30: Bullet_img = 4'd2;
//6'd14: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd14;
//6'd18,6'd19: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30: Bullet_img = 4'd1;
//6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd17,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd14;
//6'd18,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd29: Bullet_img = 4'd14;
//6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28: Bullet_img = 4'd14;
//6'd26,6'd27,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd22,6'd23: Bullet_img = 4'd13;
//6'd16,6'd18,6'd19,6'd20,6'd21,6'd24,6'd28,6'd29: Bullet_img = 4'd14;
//6'd17,6'd25,6'd26,6'd27,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd22,6'd23: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd24,6'd27,6'd28: Bullet_img = 4'd14;
//6'd25,6'd26,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd24,6'd27,6'd28,6'd29: Bullet_img = 4'd14;
//6'd25,6'd26,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd21,6'd22: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd23,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd14;
//6'd24,6'd25,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd21,6'd22: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd18,6'd19,6'd20,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd12,6'd16,6'd17,6'd24,6'd25,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd20,6'd21: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd22,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd12,6'd23,6'd24,6'd25,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd21: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd25,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd26,6'd27,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd26,6'd27,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29: Bullet_img = 4'd14;
//6'd26,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd13;
//6'd29,6'd30: Bullet_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd13;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd36: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd14;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41,6'd42: Bullet_img = 4'd2;
//6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd2;
//6'd21,6'd22,6'd23,6'd24,6'd26,6'd27: Bullet_img = 4'd4;
//6'd25: Bullet_img = 4'd12;
//6'd19: Bullet_img = 4'd13;
//6'd20,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd2;
//6'd36: Bullet_img = 4'd3;
//6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd45: Bullet_img = 4'd4;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd5;
//6'd24: Bullet_img = 4'd12;
//6'd18: Bullet_img = 4'd13;
//6'd19,6'd20,6'd44: Bullet_img = 4'd14;
//6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd2;
//6'd31,6'd32,6'd33: Bullet_img = 4'd3;
//6'd21,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd34,6'd35,6'd36: Bullet_img = 4'd5;
//6'd22,6'd23,6'd24: Bullet_img = 4'd12;
//6'd45: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20: Bullet_img = 4'd14;
//6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39: Bullet_img = 4'd2;
//6'd33: Bullet_img = 4'd3;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd32,6'd34,6'd35,6'd36: Bullet_img = 4'd5;
//6'd24,6'd25: Bullet_img = 4'd12;
//6'd21,6'd22,6'd23,6'd45: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd45: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd8;
//6'd21: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd33,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd4;
//6'd26: Bullet_img = 4'd6;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd36: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd32,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd32,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd32,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd5;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd36: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd37,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd20,6'd21: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd4;
//6'd26: Bullet_img = 4'd6;
//6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd5;
//6'd46: Bullet_img = 4'd8;
//6'd15,6'd16,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd21,6'd22,6'd23: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd45: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd24,6'd45: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd4;
//6'd19,6'd24: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd13;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd35,6'd36: Bullet_img = 4'd2;
//6'd33,6'd34: Bullet_img = 4'd3;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd32: Bullet_img = 4'd5;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35,6'd36: Bullet_img = 4'd1;
//6'd27: Bullet_img = 4'd5;
//6'd29,6'd30,6'd31: Bullet_img = 4'd13;
//6'd28,6'd32,6'd33: Bullet_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd28,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35: Bullet_img = 4'd14;
//6'd33,6'd34,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd13;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36: Bullet_img = 4'd14;
//6'd25,6'd33,6'd34,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd13;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36: Bullet_img = 4'd14;
//6'd25,6'd33,6'd34,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd25,6'd33,6'd34,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd35,6'd36,6'd37,6'd39: Bullet_img = 4'd14;
//6'd33,6'd34,6'd38,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd33,6'd34,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd32,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd25,6'd33,6'd34,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd33,6'd34,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd32,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd33,6'd34,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd30,6'd31: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd28,6'd29,6'd32,6'd33,6'd34,6'd35,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd27,6'd36,6'd37,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd31: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd32,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd26,6'd27,6'd37,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd30: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd31,6'd32: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd30: Bullet_img = 4'd13;
//6'd23,6'd24,6'd31,6'd32: Bullet_img = 4'd14;
//6'd22,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd31,6'd32,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24: Bullet_img = 4'd14;
//6'd22,6'd23: Bullet_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd35: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd14;
//6'd16,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32: Bullet_img = 4'd2;
//6'd36: Bullet_img = 4'd13;
//6'd16,6'd17,6'd22,6'd34,6'd35: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd36: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd32,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd2;
//6'd36: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26: Bullet_img = 4'd14;
//6'd24,6'd25,6'd32,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30: Bullet_img = 4'd2;
//6'd27: Bullet_img = 4'd3;
//6'd26: Bullet_img = 4'd5;
//6'd37: Bullet_img = 4'd8;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30: Bullet_img = 4'd2;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd5;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25: Bullet_img = 4'd3;
//6'd18: Bullet_img = 4'd4;
//6'd21,6'd22,6'd26,6'd27,6'd28: Bullet_img = 4'd5;
//6'd15,6'd16,6'd17,6'd19,6'd20,6'd29: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd25: Bullet_img = 4'd3;
//6'd13,6'd14,6'd17,6'd18,6'd19,6'd21,6'd22: Bullet_img = 4'd4;
//6'd20,6'd24: Bullet_img = 4'd5;
//6'd16: Bullet_img = 4'd12;
//6'd15,6'd26,6'd27,6'd28,6'd29,6'd32: Bullet_img = 4'd14;
//6'd30,6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd12;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd12;
//6'd11: Bullet_img = 4'd13;
//6'd12,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd4;
//6'd14,6'd15,6'd17,6'd18: Bullet_img = 4'd12;
//6'd16: Bullet_img = 4'd13;
//6'd11,6'd12,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10,6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd14;
//6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd31: Bullet_img = 4'd4;
//6'd20: Bullet_img = 4'd6;
//6'd15: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd32,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd31,6'd32: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd31,6'd32: Bullet_img = 4'd4;
//6'd30: Bullet_img = 4'd5;
//6'd15: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd16,6'd17,6'd18,6'd19,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd33,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd30: Bullet_img = 4'd5;
//6'd13,6'd14,6'd15: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd16,6'd17,6'd18,6'd19,6'd25,6'd26,6'd27,6'd28,6'd29,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd34,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd28,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd17,6'd18,6'd19,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd34,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd26,6'd27,6'd28,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd4;
//6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd34,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd30,6'd31,6'd33,6'd34: Bullet_img = 4'd4;
//6'd32: Bullet_img = 4'd5;
//6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd35,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28: Bullet_img = 4'd4;
//6'd45: Bullet_img = 4'd8;
//6'd15,6'd16,6'd17: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd16,6'd17,6'd18,6'd45: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd19,6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd16,6'd17,6'd18,6'd19,6'd45,6'd46: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd46: Bullet_img = 4'd4;
//6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd21,6'd22,6'd23,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27: Bullet_img = 4'd4;
//6'd28: Bullet_img = 4'd5;
//6'd26: Bullet_img = 4'd6;
//6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd22,6'd23,6'd24,6'd25,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd23: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd22,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd23,6'd24: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17,6'd24,6'd25,6'd26: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd26,6'd27: Bullet_img = 4'd13;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd2;
//6'd21,6'd22: Bullet_img = 4'd13;
//6'd20,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd1;
//6'd39: Bullet_img = 4'd2;
//6'd37,6'd38: Bullet_img = 4'd3;
//6'd21,6'd22,6'd27,6'd29,6'd30: Bullet_img = 4'd13;
//6'd23,6'd24,6'd25,6'd26,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39: Bullet_img = 4'd1;
//6'd37: Bullet_img = 4'd3;
//6'd22,6'd35: Bullet_img = 4'd4;
//6'd36: Bullet_img = 4'd5;
//6'd23,6'd26,6'd29,6'd30: Bullet_img = 4'd13;
//6'd31,6'd32,6'd33,6'd34,6'd38: Bullet_img = 4'd14;
//6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd29,6'd35,6'd36: Bullet_img = 4'd13;
//6'd37,6'd40: Bullet_img = 4'd14;
//6'd38,6'd39,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32: Bullet_img = 4'd4;
//6'd34: Bullet_img = 4'd13;
//6'd33,6'd35,6'd36,6'd37,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd38,6'd39,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd5;
//6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd33,6'd39,6'd40,6'd44,6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43,6'd44,6'd46: Bullet_img = 4'd14;
//6'd39,6'd40,6'd45,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//6'd40,6'd41,6'd47,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd31,6'd40,6'd41,6'd49,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28,6'd29,6'd30,6'd37,6'd38: Bullet_img = 4'd13;
//6'd31,6'd33,6'd34,6'd35,6'd36,6'd39,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd32,6'd40,6'd41,6'd42,6'd49,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd38,6'd39: Bullet_img = 4'd13;
//6'd31,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48: Bullet_img = 4'd14;
//6'd32,6'd41,6'd42,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd13;
//6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd40,6'd43,6'd44,6'd47,6'd48,6'd49: Bullet_img = 4'd14;
//6'd41,6'd42,6'd45,6'd46,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd38,6'd39,6'd40: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd42,6'd43,6'd44: Bullet_img = 4'd14;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd39,6'd40,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd32,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41: Bullet_img = 4'd14;
//6'd33,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd15;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd29,6'd30,6'd31,6'd32,6'd39,6'd40,6'd48,6'd49: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41: Bullet_img = 4'd14;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd40: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd41,6'd42: Bullet_img = 4'd14;
//6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd30,6'd31,6'd32,6'd33,6'd40: Bullet_img = 4'd13;
//6'd34,6'd35,6'd41,6'd42: Bullet_img = 4'd14;
//6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31,6'd32,6'd42: Bullet_img = 4'd13;
//6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd31: Bullet_img = 4'd13;
//6'd32,6'd33,6'd34: Bullet_img = 4'd14;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32: Bullet_img = 4'd13;
//6'd34,6'd35: Bullet_img = 4'd14;
//6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd13;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 12
//3'd12: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26: Bullet_img = 4'd4;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23: Bullet_img = 4'd2;
//6'd26,6'd27: Bullet_img = 4'd13;
//6'd14,6'd25: Bullet_img = 4'd14;
//6'd13: Bullet_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd27,6'd28: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd23,6'd24,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd28: Bullet_img = 4'd8;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd24,6'd25,6'd26,6'd27,6'd31: Bullet_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd2;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd2;
//6'd19: Bullet_img = 4'd3;
//6'd18: Bullet_img = 4'd14;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22: Bullet_img = 4'd2;
//6'd18,6'd19,6'd20: Bullet_img = 4'd5;
//6'd8,6'd9,6'd13,6'd14,6'd16,6'd17: Bullet_img = 4'd14;
//6'd7,6'd10,6'd11,6'd12,6'd15,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd14;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd3;
//6'd16,6'd17,6'd19,6'd20: Bullet_img = 4'd5;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd28: Bullet_img = 4'd14;
//6'd27,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19: Bullet_img = 4'd3;
//6'd15,6'd16: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd14;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16,6'd17: Bullet_img = 4'd4;
//6'd14,6'd15,6'd18: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//6'd13,6'd14: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd11,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd12;
//6'd9,6'd10,6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd14;
//6'd21,6'd28,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd27: Bullet_img = 4'd4;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd28,6'd29,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd12,6'd14,6'd27,6'd28: Bullet_img = 4'd4;
//6'd11,6'd13: Bullet_img = 4'd12;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd14;
//6'd29,6'd30,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd27,6'd28,6'd29: Bullet_img = 4'd4;
//6'd26: Bullet_img = 4'd5;
//6'd11,6'd12,6'd13: Bullet_img = 4'd12;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd30,6'd31,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd18,6'd19,6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd27: Bullet_img = 4'd5;
//6'd10: Bullet_img = 4'd12;
//6'd11,6'd12: Bullet_img = 4'd13;
//6'd7,6'd8,6'd13,6'd14,6'd15,6'd16,6'd17,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd31,6'd32,6'd37,6'd38,6'd39,6'd40,6'd41,6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd6;
//6'd10,6'd11,6'd12,6'd44: Bullet_img = 4'd13;
//6'd7,6'd8,6'd9,6'd13,6'd14,6'd15,6'd16,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd32,6'd33,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd21,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd4;
//6'd6,6'd7,6'd11,6'd44,6'd45: Bullet_img = 4'd13;
//6'd8,6'd9,6'd10,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd22,6'd23,6'd24,6'd25,6'd26,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd25,6'd26,6'd28,6'd45: Bullet_img = 4'd4;
//6'd30: Bullet_img = 4'd5;
//6'd12: Bullet_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd13,6'd14,6'd15,6'd16,6'd22,6'd23,6'd24,6'd27,6'd29,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd14,6'd15,6'd16,6'd17,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd25,6'd26: Bullet_img = 4'd4;
//6'd12,6'd13: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd14,6'd15,6'd16,6'd17,6'd20,6'd21,6'd22,6'd23,6'd24,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd14: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd13;
//6'd10,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27: Bullet_img = 4'd4;
//6'd12,6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd13,6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd4;
//6'd14,6'd15,6'd16,6'd17,6'd18: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd19,6'd20,6'd21,6'd22,6'd23,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd4;
//6'd30: Bullet_img = 4'd5;
//6'd15,6'd16,6'd17,6'd18,6'd19: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd29: Bullet_img = 4'd5;
//6'd28: Bullet_img = 4'd6;
//6'd16,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd21,6'd22,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43: Bullet_img = 4'd2;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: Bullet_img = 4'd13;
//6'd13,6'd14,6'd15,6'd16,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd1;
//6'd42,6'd43: Bullet_img = 4'd2;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd14;
//6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43: Bullet_img = 4'd1;
//6'd41,6'd42: Bullet_img = 4'd3;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd44,6'd47,6'd51: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd3;
//6'd40: Bullet_img = 4'd5;
//6'd20,6'd21,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd13;
//6'd16,6'd17,6'd18,6'd19,6'd22,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd42,6'd45,6'd46,6'd50: Bullet_img = 4'd14;
//6'd43,6'd44,6'd47,6'd48,6'd49,6'd51,6'd52,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40: Bullet_img = 4'd4;
//6'd24,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd41,6'd45,6'd46,6'd47,6'd48,6'd49,6'd51: Bullet_img = 4'd14;
//6'd42,6'd43,6'd44,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd38,6'd39: Bullet_img = 4'd4;
//6'd28,6'd34,6'd40: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd43,6'd44,6'd45,6'd55,6'd56,6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd37,6'd38: Bullet_img = 4'd4;
//6'd36: Bullet_img = 4'd12;
//6'd32,6'd33,6'd34,6'd35,6'd39: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd44,6'd45,6'd46,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37: Bullet_img = 4'd4;
//6'd21,6'd22,6'd31,6'd34,6'd59: Bullet_img = 4'd13;
//6'd20,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd38,6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55: Bullet_img = 4'd14;
//6'd39,6'd45,6'd46,6'd47,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd21,6'd22,6'd26,6'd27,6'd28,6'd29,6'd38,6'd58,6'd59: Bullet_img = 4'd13;
//6'd25,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd49,6'd50,6'd51,6'd54: Bullet_img = 4'd14;
//6'd39,6'd46,6'd47,6'd48,6'd52,6'd53,6'd55,6'd56,6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28: Bullet_img = 4'd4;
//6'd44,6'd45,6'd57,6'd58: Bullet_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd46,6'd50,6'd51: Bullet_img = 4'd14;
//6'd47,6'd48,6'd49,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd44,6'd45,6'd46,6'd56,6'd57: Bullet_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd47,6'd50,6'd51: Bullet_img = 4'd14;
//6'd48,6'd49,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd45,6'd46,6'd47: Bullet_img = 4'd13;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd48,6'd49,6'd50: Bullet_img = 4'd14;
//6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd46,6'd47,6'd48: Bullet_img = 4'd13;
//6'd38,6'd41,6'd42,6'd43,6'd44,6'd45,6'd49: Bullet_img = 4'd14;
//6'd39,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36,6'd37,6'd38,6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//6'd39,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd50: Bullet_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd39,6'd49: Bullet_img = 4'd13;
//6'd38,6'd40,6'd41,6'd43,6'd44,6'd45,6'd46,6'd47,6'd50,6'd51: Bullet_img = 4'd14;
//6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd37,6'd38,6'd39,6'd40,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd13;
//6'd41,6'd43,6'd44,6'd46: Bullet_img = 4'd14;
//6'd42,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd13;
//6'd42,6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd13;
//6'd43,6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd13;
//6'd44,6'd45,6'd46: Bullet_img = 4'd14;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd41,6'd42: Bullet_img = 4'd13;
//6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd42,6'd46: Bullet_img = 4'd13;
//6'd43,6'd44,6'd45: Bullet_img = 4'd14;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43,6'd45,6'd46: Bullet_img = 4'd13;
//6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd13;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 13
//3'd13: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17: Bullet_img = 4'd4;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18,6'd19,6'd20: Bullet_img = 4'd13;
//6'd17: Bullet_img = 4'd14;
//6'd21: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14: Bullet_img = 4'd2;
//6'd20,6'd21: Bullet_img = 4'd8;
//6'd24,6'd25: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15: Bullet_img = 4'd2;
//6'd16,6'd17,6'd18,6'd19,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14: Bullet_img = 4'd2;
//6'd11,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//6'd7: Bullet_img = 4'd14;
//6'd6,6'd8,6'd9,6'd10,6'd11,6'd12,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd2;
//6'd39: Bullet_img = 4'd8;
//6'd19,6'd20,6'd21,6'd22,6'd23: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd17,6'd18,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15: Bullet_img = 4'd5;
//6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd40: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15: Bullet_img = 4'd5;
//6'd41: Bullet_img = 4'd13;
//6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd14;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd43: Bullet_img = 4'd4;
//6'd12,6'd13,6'd14,6'd15: Bullet_img = 4'd5;
//6'd42: Bullet_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd14;
//6'd4,6'd5,6'd6,6'd7,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14: Bullet_img = 4'd3;
//6'd12: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd11,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd24,6'd25,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd3;
//6'd23,6'd24,6'd25: Bullet_img = 4'd4;
//6'd12,6'd14: Bullet_img = 4'd5;
//6'd4,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd14;
//6'd3,6'd5,6'd26,6'd27,6'd28,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd5;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd14,6'd15,6'd16,6'd17,6'd19,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd3,6'd18,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd12,6'd13,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd4;
//6'd11,6'd24,6'd25: Bullet_img = 4'd5;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd11,6'd12,6'd13,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd4;
//6'd10: Bullet_img = 4'd5;
//6'd5,6'd6,6'd7,6'd8,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12,6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd28: Bullet_img = 4'd5;
//6'd5,6'd6,6'd7,6'd8,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36: Bullet_img = 4'd14;
//6'd37,6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd4;
//6'd8: Bullet_img = 4'd12;
//default: Bullet_img = 4'd14;
//6'd38,6'd39,6'd40,6'd41: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd8,6'd9,6'd10,6'd17,6'd18,6'd19,6'd24,6'd25,6'd26: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd12;
//6'd7,6'd12,6'd13,6'd14,6'd15,6'd16,6'd20,6'd21,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd7,6'd8,6'd17,6'd18,6'd19,6'd20,6'd21,6'd24,6'd25,6'd26: Bullet_img = 4'd4;
//6'd16: Bullet_img = 4'd6;
//6'd9,6'd10,6'd11: Bullet_img = 4'd12;
//6'd12,6'd13,6'd14,6'd15,6'd22,6'd23,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd6,6'd7,6'd8,6'd17,6'd18,6'd19,6'd20,6'd24,6'd25,6'd26: Bullet_img = 4'd4;
//6'd9,6'd11: Bullet_img = 4'd12;
//6'd10: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd47,6'd48,6'd50,6'd63,6'd64: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd1;
//6'd45: Bullet_img = 4'd2;
//6'd6,6'd7,6'd8,6'd17,6'd18,6'd19,6'd20: Bullet_img = 4'd4;
//6'd9: Bullet_img = 4'd12;
//6'd10,6'd11,6'd62: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd40,6'd41,6'd42,6'd43,6'd44,6'd49,6'd51,6'd52,6'd58,6'd59,6'd60,6'd61: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd63,6'd64: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd1;
//6'd44: Bullet_img = 4'd3;
//6'd8,6'd9,6'd18,6'd19,6'd27,6'd28: Bullet_img = 4'd4;
//6'd10,6'd11,6'd62: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd41,6'd42,6'd43,6'd46,6'd48,6'd50,6'd59,6'd60,6'd61: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd45: Bullet_img = 4'd1;
//6'd44: Bullet_img = 4'd3;
//6'd19,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd6,6'd11,6'd12,6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd42,6'd43,6'd46,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd32,6'd43,6'd44: Bullet_img = 4'd5;
//6'd7,6'd13,6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd46,6'd47,6'd48,6'd49,6'd56,6'd57,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd59,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd43: Bullet_img = 4'd4;
//6'd31: Bullet_img = 4'd5;
//6'd30: Bullet_img = 4'd6;
//6'd13,6'd14,6'd15,6'd60: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd56,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd26,6'd27,6'd28,6'd29,6'd43: Bullet_img = 4'd4;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd44: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd42: Bullet_img = 4'd4;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd43: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd42: Bullet_img = 4'd4;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd32,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd40,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd4;
//6'd42,6'd43: Bullet_img = 4'd5;
//default: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd36,6'd37,6'd45,6'd46,6'd47,6'd48,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//6'd44: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd40,6'd42,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd41: Bullet_img = 4'd4;
//default: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd33,6'd34,6'd35,6'd36,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd56,6'd57: Bullet_img = 4'd14;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd22,6'd23,6'd24,6'd25,6'd27,6'd28,6'd29,6'd30,6'd36,6'd44,6'd54,6'd58: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd26,6'd31,6'd32,6'd33,6'd34,6'd35,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd56,6'd57: Bullet_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd25,6'd36,6'd43,6'd56: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd44,6'd45: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd43: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd45,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34: Bullet_img = 4'd4;
//6'd32,6'd33,6'd44: Bullet_img = 4'd13;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd45,6'd46,6'd47,6'd48,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd49,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd29,6'd43,6'd44,6'd46,6'd47: Bullet_img = 4'd13;
//6'd24,6'd25,6'd26,6'd45,6'd48,6'd49,6'd50,6'd51,6'd52,6'd54: Bullet_img = 4'd14;
//6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd27,6'd28,6'd46,6'd47,6'd48,6'd49: Bullet_img = 4'd13;
//6'd45,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51: Bullet_img = 4'd13;
//6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd55: Bullet_img = 4'd13;
//6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd49,6'd50,6'd51,6'd55: Bullet_img = 4'd13;
//6'd52: Bullet_img = 4'd14;
//6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd52,6'd53,6'd54: Bullet_img = 4'd13;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 14
//3'd14: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34: Bullet_img = 4'd8;
//6'd15,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd36: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd39: Bullet_img = 4'd4;
//6'd15: Bullet_img = 4'd8;
//6'd12,6'd13,6'd14,6'd37,6'd38: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11: Bullet_img = 4'd14;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd39: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd9,6'd10: Bullet_img = 4'd2;
//6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd40,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd9,6'd10: Bullet_img = 4'd2;
//6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd2;
//6'd61: Bullet_img = 4'd13;
//6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd52,6'd53,6'd54,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd7,6'd8,6'd9,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd51,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd41,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd7,6'd8,6'd9,6'd14,6'd15,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd51,6'd52,6'd59,6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13: Bullet_img = 4'd2;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd44,6'd47,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd1;
//6'd10,6'd45: Bullet_img = 4'd2;
//6'd11: Bullet_img = 4'd3;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29: Bullet_img = 4'd4;
//6'd12,6'd13: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd40,6'd41,6'd42,6'd43,6'd48,6'd57: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd1;
//6'd45: Bullet_img = 4'd2;
//6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd4;
//6'd11,6'd12,6'd13: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd41,6'd42,6'd43,6'd44,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd46: Bullet_img = 4'd1;
//6'd45: Bullet_img = 4'd3;
//6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd11,6'd12,6'd13,6'd23,6'd24,6'd28: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd41,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd2,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd12,6'd13,6'd45: Bullet_img = 4'd3;
//6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd17,6'd42,6'd43,6'd44,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd3;
//6'd11,6'd13,6'd45: Bullet_img = 4'd5;
//6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd12: Bullet_img = 4'd3;
//6'd13,6'd25,6'd26,6'd27,6'd45: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd5;
//6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd2,6'd58,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd12,6'd13,6'd25,6'd26,6'd27,6'd45: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd5;
//6'd46,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd59,6'd60: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5,6'd6: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//6'd1,6'd2,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd12,6'd13,6'd25,6'd26,6'd27,6'd45: Bullet_img = 4'd4;
//6'd11: Bullet_img = 4'd5;
//6'd46: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd4,6'd5: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//6'd1,6'd2,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd12,6'd13,6'd18,6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd45: Bullet_img = 4'd4;
//6'd11,6'd34: Bullet_img = 4'd5;
//default: Bullet_img = 4'd14;
//6'd3,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//6'd1,6'd2,6'd44,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd33,6'd45: Bullet_img = 4'd4;
//6'd34,6'd46: Bullet_img = 4'd5;
//6'd47: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd3,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd44,6'd46,6'd47,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd10,6'd11,6'd12,6'd13,6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32,6'd45: Bullet_img = 4'd4;
//6'd18,6'd33: Bullet_img = 4'd6;
//6'd42,6'd43,6'd48: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd44,6'd45,6'd46,6'd47,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd11,6'd12,6'd19,6'd20,6'd21,6'd22,6'd29,6'd30,6'd31,6'd32: Bullet_img = 4'd4;
//6'd10,6'd13: Bullet_img = 4'd12;
//6'd42,6'd43,6'd48: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd10,6'd21,6'd22,6'd29,6'd30,6'd31: Bullet_img = 4'd4;
//6'd11,6'd12,6'd13: Bullet_img = 4'd12;
//6'd36,6'd37,6'd38,6'd39,6'd41,6'd48,6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//endcase
//end
//6'd41: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd12;
//6'd13,6'd14,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//endcase
//end
//6'd42: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd42,6'd43,6'd44,6'd45,6'd46,6'd47,6'd48,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd12;
//6'd13,6'd14,6'd33,6'd34,6'd35,6'd36,6'd37,6'd41,6'd49,6'd50,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd61: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd60: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd4;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd51,6'd52,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd36,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd40: Bullet_img = 4'd4;
//6'd10,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd38,6'd39: Bullet_img = 4'd13;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd11,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd38: Bullet_img = 4'd13;
//6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd36: Bullet_img = 4'd13;
//6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd34,6'd35: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//// Bullet_type_2 15
//3'd15: begin
//case(y)
//6'd0: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd1: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd2: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd3: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd4: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd5: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd6: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd7: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd8: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd9: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd10: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd11: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd55: Bullet_img = 4'd13;
//endcase
//end
//6'd12: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd55: Bullet_img = 4'd13;
//6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd55: Bullet_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd56: Bullet_img = 4'd13;
//6'd53: Bullet_img = 4'd14;
//6'd49,6'd50,6'd51,6'd52,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd56: Bullet_img = 4'd13;
//6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd14;
//6'd48,6'd49,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd33: Bullet_img = 4'd4;
//6'd32: Bullet_img = 4'd13;
//6'd48,6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd30,6'd47,6'd53,6'd54,6'd55: Bullet_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd28: Bullet_img = 4'd8;
//6'd31,6'd32: Bullet_img = 4'd13;
//6'd49,6'd50,6'd51,6'd52: Bullet_img = 4'd14;
//6'd27,6'd34,6'd47,6'd48,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd33,6'd47: Bullet_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd14;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd46: Bullet_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd59: Bullet_img = 4'd13;
//6'd46,6'd47,6'd48,6'd49,6'd50,6'd54,6'd57,6'd58: Bullet_img = 4'd14;
//6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd46,6'd47,6'd48,6'd54,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd14;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd45,6'd49,6'd50,6'd51,6'd52,6'd53: Bullet_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd38,6'd39,6'd40,6'd41,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd43: Bullet_img = 4'd1;
//6'd42: Bullet_img = 4'd2;
//6'd54,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd13;
//6'd45,6'd46,6'd52,6'd53: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd1;
//6'd43: Bullet_img = 4'd2;
//6'd52,6'd53,6'd54,6'd55,6'd56: Bullet_img = 4'd13;
//6'd28,6'd29,6'd49,6'd50,6'd51: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd12,6'd13,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd43: Bullet_img = 4'd3;
//6'd51,6'd52,6'd53,6'd54: Bullet_img = 4'd13;
//6'd26,6'd27,6'd28,6'd29,6'd30,6'd37,6'd44,6'd47,6'd48,6'd49,6'd50,6'd55,6'd56: Bullet_img = 4'd14;
//default: Bullet_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd12,6'd57,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd43,6'd44: Bullet_img = 4'd3;
//6'd11: Bullet_img = 4'd8;
//6'd51: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd39,6'd40,6'd41,6'd42,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd11,6'd12,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd44: Bullet_img = 4'd5;
//6'd8,6'd9,6'd10,6'd45: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd41,6'd57,6'd58: Bullet_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd9,6'd10,6'd60,6'd63,6'd64: Bullet_img = 4'd0;
//6'd7,6'd44: Bullet_img = 4'd4;
//6'd45,6'd62: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd27: Bullet_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd9,6'd63,6'd64: Bullet_img = 4'd0;
//6'd27,6'd45: Bullet_img = 4'd4;
//6'd46,6'd62: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd24,6'd25,6'd26: Bullet_img = 4'd15;
//endcase
//end
//6'd30: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd63,6'd64: Bullet_img = 4'd0;
//6'd24,6'd25,6'd26,6'd27,6'd45: Bullet_img = 4'd4;
//6'd58,6'd62: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd22,6'd23,6'd47,6'd55,6'd61: Bullet_img = 4'd15;
//endcase
//end
//6'd31: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd48,6'd63,6'd64: Bullet_img = 4'd0;
//6'd7,6'd8: Bullet_img = 4'd2;
//6'd22,6'd23,6'd24,6'd25,6'd26,6'd45,6'd46: Bullet_img = 4'd4;
//6'd27,6'd47: Bullet_img = 4'd5;
//6'd49,6'd56,6'd57,6'd58,6'd59,6'd61,6'd62: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd21,6'd51,6'd52: Bullet_img = 4'd15;
//endcase
//end
//6'd32: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd45,6'd47,6'd48,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd2;
//6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd46: Bullet_img = 4'd4;
//6'd49,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd11,6'd12,6'd13,6'd14,6'd50: Bullet_img = 4'd15;
//endcase
//end
//6'd33: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd45,6'd46,6'd47,6'd48,6'd49,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd2;
//6'd25,6'd26,6'd27: Bullet_img = 4'd4;
//6'd23,6'd24: Bullet_img = 4'd5;
//6'd43,6'd44,6'd50,6'd51,6'd52,6'd54,6'd55,6'd56,6'd57,6'd58: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd13,6'd14: Bullet_img = 4'd15;
//endcase
//end
//6'd34: begin
//case(x)
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd46,6'd47,6'd48,6'd49,6'd50,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11,6'd12: Bullet_img = 4'd2;
//6'd43,6'd44,6'd45,6'd51,6'd52,6'd54,6'd55,6'd56: Bullet_img = 4'd13;
//default: Bullet_img = 4'd14;
//6'd7,6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd35: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd9,6'd10,6'd11: Bullet_img = 4'd2;
//6'd25,6'd26,6'd27,6'd28,6'd33,6'd34: Bullet_img = 4'd4;
//6'd12,6'd13,6'd35: Bullet_img = 4'd5;
//6'd51: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd29,6'd30,6'd31,6'd32,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd6,6'd7,6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd36: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd10: Bullet_img = 4'd2;
//6'd11: Bullet_img = 4'd3;
//6'd26,6'd27,6'd28,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd4;
//6'd12,6'd13: Bullet_img = 4'd5;
//6'd41,6'd43: Bullet_img = 4'd13;
//6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd29,6'd30,6'd36,6'd37,6'd38,6'd39,6'd40,6'd42: Bullet_img = 4'd14;
//6'd6,6'd7,6'd8,6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd37: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd26,6'd27,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd11,6'd12,6'd13: Bullet_img = 4'd5;
//6'd35: Bullet_img = 4'd6;
//6'd39,6'd40,6'd41,6'd44: Bullet_img = 4'd13;
//6'd10,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd28,6'd29,6'd30,6'd36,6'd37,6'd38,6'd42,6'd43: Bullet_img = 4'd14;
//6'd6,6'd7,6'd8,6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd38: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14: Bullet_img = 4'd3;
//6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd5;
//6'd39,6'd40: Bullet_img = 4'd13;
//6'd11,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd35,6'd36,6'd37,6'd38,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd15;
//endcase
//end
//6'd39: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13: Bullet_img = 4'd3;
//6'd24,6'd31,6'd32,6'd33,6'd34: Bullet_img = 4'd4;
//6'd12,6'd14: Bullet_img = 4'd5;
//6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd13;
//6'd4,6'd11,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd35,6'd36,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8,6'd9,6'd10: Bullet_img = 4'd15;
//endcase
//end
//6'd40: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14: Bullet_img = 4'd3;
//6'd15,6'd21,6'd22,6'd23,6'd24,6'd32,6'd33: Bullet_img = 4'd4;
//6'd12: Bullet_img = 4'd5;
//6'd36,6'd37,6'd38,6'd39,6'd44: Bullet_img = 4'd13;
//6'd10,6'd11,6'd16,6'd17,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd34,6'd35,6'd40,6'd41,6'd42,6'd43: Bullet_img = 4'd14;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9: Bullet_img = 4'd15;
//endcase
//end
//6'd41: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd44: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd5;
//6'd37,6'd38,6'd39,6'd42,6'd43: Bullet_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd16,6'd17,6'd18,6'd19,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd40,6'd41: Bullet_img = 4'd14;
//6'd4,6'd5,6'd6,6'd7: Bullet_img = 4'd15;
//endcase
//end
//6'd42: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd21,6'd22,6'd23,6'd24,6'd25: Bullet_img = 4'd4;
//6'd13: Bullet_img = 4'd5;
//6'd35,6'd36,6'd37,6'd38,6'd42,6'd43: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd16,6'd17,6'd18,6'd19,6'd20,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd39,6'd40,6'd41: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd43: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16,6'd22,6'd23,6'd24,6'd25,6'd26: Bullet_img = 4'd4;
//6'd14: Bullet_img = 4'd5;
//6'd21: Bullet_img = 4'd6;
//6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd38,6'd39,6'd40,6'd41,6'd42: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd44: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd32,6'd33,6'd34,6'd35,6'd36,6'd41: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd13,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd5,6'd6,6'd7,6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd45: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd13,6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd12;
//6'd30,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd41: Bullet_img = 4'd13;
//6'd9,6'd10,6'd11,6'd12,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd37,6'd38,6'd39,6'd40: Bullet_img = 4'd14;
//6'd6,6'd7,6'd8: Bullet_img = 4'd15;
//endcase
//end
//6'd46: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd12;
//6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd40,6'd41: Bullet_img = 4'd13;
//6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd6: Bullet_img = 4'd15;
//endcase
//end
//6'd47: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd12;
//6'd17,6'd18,6'd19,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd40: Bullet_img = 4'd13;
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd20,6'd21,6'd22,6'd23,6'd24,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39: Bullet_img = 4'd14;
//6'd7: Bullet_img = 4'd15;
//endcase
//end
//6'd48: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15,6'd16: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd12;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd13;
//6'd10,6'd11,6'd12,6'd13,6'd14,6'd31,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37: Bullet_img = 4'd14;
//endcase
//end
//6'd49: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16: Bullet_img = 4'd4;
//6'd17: Bullet_img = 4'd12;
//6'd18,6'd19,6'd24,6'd25,6'd26,6'd27: Bullet_img = 4'd13;
//6'd12,6'd20,6'd21,6'd22,6'd23,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd35: Bullet_img = 4'd14;
//endcase
//end
//6'd50: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd14,6'd15,6'd16,6'd17: Bullet_img = 4'd4;
//6'd24,6'd25: Bullet_img = 4'd13;
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd26,6'd27,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33: Bullet_img = 4'd14;
//endcase
//end
//6'd51: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd15: Bullet_img = 4'd4;
//6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30: Bullet_img = 4'd14;
//endcase
//end
//6'd52: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd16: Bullet_img = 4'd13;
//6'd17,6'd18,6'd19,6'd20,6'd22,6'd23,6'd24,6'd25,6'd26,6'd27,6'd28: Bullet_img = 4'd14;
//endcase
//end
//6'd53: begin
//case(x)
//default: Bullet_img = 4'd0;
//6'd18: Bullet_img = 4'd13;
//6'd24,6'd25: Bullet_img = 4'd14;
//endcase
//end
//6'd54: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd55: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd56: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd57: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd58: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd59: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd60: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd61: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd62: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//6'd63: begin
//case(x)
//default: Bullet_img = 4'd0;
//endcase
//end
//endcase
//end
//endcase
//
//end
//endcase
end
endfunction
function [3:0] GUI_img(input [6:0] x, input [6:0] y, input [3:0] e_type);
begin
//case(e_type)
//// Element_type 0
//3'd0: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 1
//3'd1: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 2
//3'd2: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 3
//3'd3: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 4
//3'd4: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 5
//3'd5: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 6
//3'd6: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd18,6'd19,6'd20,6'd21,6'd22,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 7
//3'd7: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 8
//3'd8: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 9
//3'd9: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//default: GUI_img = 4'd12;
//6'd1,6'd2,6'd3,6'd4,6'd5,6'd6,6'd7,6'd23,6'd24: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd29: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 10
//3'd10: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd21,6'd22: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85,6'd86,6'd87,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85,6'd86,6'd87,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85,6'd86,6'd87,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85,6'd86,6'd87,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd83,6'd84,6'd85,6'd86,6'd87,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd93,6'd94,6'd95,6'd96,6'd97,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd93,6'd94,6'd95,6'd96,6'd97,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd93,6'd94,6'd95,6'd96,6'd97,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd93,6'd94,6'd95,6'd96,6'd97,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd78,6'd79,6'd80,6'd81,6'd82,6'd93,6'd94,6'd95,6'd96,6'd97,6'd103,6'd104,6'd105,6'd106,6'd107,6'd108,6'd109,6'd110,6'd111,6'd112: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd18,6'd19,6'd20,6'd21,6'd22,6'd28,6'd29,6'd30,6'd31,6'd32,6'd48,6'd49,6'd50,6'd51,6'd52,6'd63,6'd64,6'd65,6'd66,6'd67,6'd73,6'd74,6'd75,6'd76,6'd77,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd3,6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd33,6'd34,6'd35,6'd36,6'd37,6'd38,6'd39,6'd40,6'd41,6'd42,6'd53,6'd54,6'd55,6'd56,6'd57,6'd58,6'd59,6'd60,6'd61,6'd62,6'd73,6'd74,6'd75,6'd76,6'd77,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105,6'd106,6'd107: GUI_img = 4'd12;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//// Element_type 11
//3'd11: begin
//case(y)
//6'd0: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd1: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd2: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20: GUI_img = 4'd12;
//6'd3,6'd17: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd3: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20: GUI_img = 4'd12;
//6'd3,6'd17: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd4: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20: GUI_img = 4'd12;
//6'd3,6'd17: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd5: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20: GUI_img = 4'd12;
//6'd3,6'd17: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd6: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//6'd3,6'd17,6'd55,6'd58,6'd92: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd7: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//6'd3,6'd17,6'd55,6'd58,6'd92: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd8: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102: GUI_img = 4'd12;
//6'd3,6'd17,6'd55,6'd58,6'd92: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd9: begin
//case(x)
//6'd4,6'd5,6'd6,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95: GUI_img = 4'd12;
//6'd3,6'd11,6'd12,6'd13,6'd17,6'd24,6'd31,6'd38,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd96,6'd97,6'd98,6'd99,6'd100,6'd101,6'd102,6'd103,6'd104,6'd105: GUI_img = 4'd13;
//6'd10,6'd106: GUI_img = 4'd14;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd10: begin
//case(x)
//6'd4,6'd5,6'd6,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd3,6'd10,6'd17,6'd24,6'd31,6'd38,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd11: begin
//case(x)
//6'd4,6'd5,6'd6,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd3,6'd10,6'd17,6'd24,6'd31,6'd38,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd12: begin
//case(x)
//6'd4,6'd5,6'd6,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd32,6'd33,6'd34,6'd35,6'd36,6'd37,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd3,6'd10,6'd17,6'd24,6'd31,6'd38,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd13: begin
//case(x)
//6'd4,6'd5,6'd6,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd3,6'd10,6'd17,6'd24,6'd31,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd14: begin
//case(x)
//6'd4,6'd5,6'd6,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd3,6'd10,6'd17,6'd24,6'd31,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd15: begin
//case(x)
//6'd4,6'd5,6'd6,6'd11,6'd12,6'd13,6'd18,6'd19,6'd20,6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd42,6'd43,6'd44,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd69,6'd70,6'd71,6'd76,6'd77,6'd78,6'd86,6'd87,6'd88,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd3,6'd10,6'd17,6'd24,6'd31,6'd41,6'd55,6'd58,6'd72,6'd75,6'd89,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd16: begin
//case(x)
//6'd25,6'd26,6'd27,6'd28,6'd29,6'd30,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd4,6'd5,6'd6,6'd7,6'd8,6'd9,6'd10,6'd11,6'd12,6'd13,6'd14,6'd15,6'd16,6'd17,6'd18,6'd19,6'd20,6'd24,6'd31,6'd55,6'd58,6'd92,6'd106: GUI_img = 4'd13;
//6'd3: GUI_img = 4'd14;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd17: begin
//case(x)
//6'd7,6'd8,6'd9,6'd14,6'd15,6'd16,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd10,6'd17,6'd55,6'd58,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd18: begin
//case(x)
//6'd7,6'd8,6'd9,6'd14,6'd15,6'd16,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd10,6'd17,6'd55,6'd58,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd19: begin
//case(x)
//6'd7,6'd8,6'd9,6'd14,6'd15,6'd16,6'd28,6'd29,6'd30,6'd31,6'd32,6'd33,6'd34,6'd45,6'd46,6'd47,6'd48,6'd49,6'd50,6'd51,6'd52,6'd53,6'd54,6'd59,6'd60,6'd61,6'd62,6'd63,6'd64,6'd65,6'd66,6'd67,6'd68,6'd79,6'd80,6'd81,6'd82,6'd83,6'd84,6'd85,6'd93,6'd94,6'd95,6'd103,6'd104,6'd105: GUI_img = 4'd12;
//6'd10,6'd17,6'd55,6'd58,6'd92,6'd106: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd20: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd21: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd22: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd23: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd24: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd25: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd26: begin
//case(x)
//6'd59,6'd60,6'd61: GUI_img = 4'd12;
//6'd58: GUI_img = 4'd13;
//default: GUI_img = 4'd15;
//endcase
//end
//6'd27: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//6'd28: begin
//case(x)
//default: GUI_img = 4'd15;
//endcase
//end
//endcase
//end
//endcase

end
endfunction
endmodule
