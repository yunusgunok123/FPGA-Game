module GUI_init (
		output reg[3:0] Number0 [0:23][0:29],
		output reg[3:0] Number1 [0:23][0:29],
		output reg[3:0] Number2 [0:23][0:29],
		output reg[3:0] Number3 [0:23][0:29],
		output reg[3:0] Number4 [0:23][0:29],
		output reg[3:0] Number5 [0:23][0:29],
		output reg[3:0] Number6 [0:23][0:29],
		output reg[3:0] Number7 [0:23][0:29],
		output reg[3:0] Number8 [0:23][0:29],
		output reg[3:0] Number9 [0:23][0:29],
		output reg[3:0] S_A [0:114][0:28], // Score article image
		output reg[3:0] W_A [0:107][0:28] // Weapon article image
);

initial begin

// Storing the pixel color information of Pictures of numbers for Score

//Number 0
    Number0[0][0] = 4'hF;
    Number0[1][0] = 4'hF;
    Number0[2][0] = 4'hF;
    Number0[3][0] = 4'hF;
    Number0[4][0] = 4'hF;
    Number0[5][0] = 4'hF;
    Number0[6][0] = 4'hF;
    Number0[7][0] = 4'hF;
    Number0[8][0] = 4'hF;
    Number0[9][0] = 4'hF;
    Number0[10][0] = 4'hF;
    Number0[11][0] = 4'hF;
    Number0[12][0] = 4'hF;
    Number0[13][0] = 4'hF;
    Number0[14][0] = 4'hF;
    Number0[15][0] = 4'hF;
    Number0[16][0] = 4'hF;
    Number0[17][0] = 4'hF;
    Number0[18][0] = 4'hF;
    Number0[19][0] = 4'hF;
    Number0[20][0] = 4'hF;
    Number0[21][0] = 4'hF;
    Number0[22][0] = 4'hF;
    Number0[23][0] = 4'hF;
    Number0[0][1] = 4'hF;
    Number0[1][1] = 4'hF;
    Number0[2][1] = 4'hF;
    Number0[3][1] = 4'hF;
    Number0[4][1] = 4'hF;
    Number0[5][1] = 4'hF;
    Number0[6][1] = 4'hF;
    Number0[7][1] = 4'hF;
    Number0[8][1] = 4'hF;
    Number0[9][1] = 4'hF;
    Number0[10][1] = 4'hF;
    Number0[11][1] = 4'hF;
    Number0[12][1] = 4'hF;
    Number0[13][1] = 4'hF;
    Number0[14][1] = 4'hF;
    Number0[15][1] = 4'hF;
    Number0[16][1] = 4'hF;
    Number0[17][1] = 4'hF;
    Number0[18][1] = 4'hF;
    Number0[19][1] = 4'hF;
    Number0[20][1] = 4'hF;
    Number0[21][1] = 4'hF;
    Number0[22][1] = 4'hF;
    Number0[23][1] = 4'hF;
    Number0[0][2] = 4'hF;
    Number0[1][2] = 4'hF;
    Number0[2][2] = 4'hF;
    Number0[3][2] = 4'hF;
    Number0[4][2] = 4'hF;
    Number0[5][2] = 4'hF;
    Number0[6][2] = 4'hF;
    Number0[7][2] = 4'hF;
    Number0[8][2] = 4'hF;
    Number0[9][2] = 4'hF;
    Number0[10][2] = 4'hF;
    Number0[11][2] = 4'hF;
    Number0[12][2] = 4'hF;
    Number0[13][2] = 4'hF;
    Number0[14][2] = 4'hF;
    Number0[15][2] = 4'hF;
    Number0[16][2] = 4'hF;
    Number0[17][2] = 4'hF;
    Number0[18][2] = 4'hF;
    Number0[19][2] = 4'hF;
    Number0[20][2] = 4'hF;
    Number0[21][2] = 4'hF;
    Number0[22][2] = 4'hF;
    Number0[23][2] = 4'hF;
    Number0[0][3] = 4'hF;
    Number0[1][3] = 4'hF;
    Number0[2][3] = 4'hF;
    Number0[3][3] = 4'hF;
    Number0[4][3] = 4'hF;
    Number0[5][3] = 4'hF;
    Number0[6][3] = 4'hF;
    Number0[7][3] = 4'hC;
    Number0[8][3] = 4'hC;
    Number0[9][3] = 4'hC;
    Number0[10][3] = 4'hC;
    Number0[11][3] = 4'hC;
    Number0[12][3] = 4'hC;
    Number0[13][3] = 4'hC;
    Number0[14][3] = 4'hC;
    Number0[15][3] = 4'hC;
    Number0[16][3] = 4'hC;
    Number0[17][3] = 4'hF;
    Number0[18][3] = 4'hF;
    Number0[19][3] = 4'hF;
    Number0[20][3] = 4'hF;
    Number0[21][3] = 4'hF;
    Number0[22][3] = 4'hF;
    Number0[23][3] = 4'hF;
    Number0[0][4] = 4'hF;
    Number0[1][4] = 4'hF;
    Number0[2][4] = 4'hF;
    Number0[3][4] = 4'hF;
    Number0[4][4] = 4'hF;
    Number0[5][4] = 4'hF;
    Number0[6][4] = 4'hF;
    Number0[7][4] = 4'hC;
    Number0[8][4] = 4'hC;
    Number0[9][4] = 4'hC;
    Number0[10][4] = 4'hC;
    Number0[11][4] = 4'hC;
    Number0[12][4] = 4'hC;
    Number0[13][4] = 4'hC;
    Number0[14][4] = 4'hC;
    Number0[15][4] = 4'hC;
    Number0[16][4] = 4'hC;
    Number0[17][4] = 4'hF;
    Number0[18][4] = 4'hF;
    Number0[19][4] = 4'hF;
    Number0[20][4] = 4'hF;
    Number0[21][4] = 4'hF;
    Number0[22][4] = 4'hF;
    Number0[23][4] = 4'hF;
    Number0[0][5] = 4'hF;
    Number0[1][5] = 4'hF;
    Number0[2][5] = 4'hF;
    Number0[3][5] = 4'hF;
    Number0[4][5] = 4'hF;
    Number0[5][5] = 4'hF;
    Number0[6][5] = 4'hF;
    Number0[7][5] = 4'hC;
    Number0[8][5] = 4'hC;
    Number0[9][5] = 4'hC;
    Number0[10][5] = 4'hC;
    Number0[11][5] = 4'hC;
    Number0[12][5] = 4'hC;
    Number0[13][5] = 4'hC;
    Number0[14][5] = 4'hC;
    Number0[15][5] = 4'hC;
    Number0[16][5] = 4'hC;
    Number0[17][5] = 4'hF;
    Number0[18][5] = 4'hF;
    Number0[19][5] = 4'hF;
    Number0[20][5] = 4'hF;
    Number0[21][5] = 4'hF;
    Number0[22][5] = 4'hF;
    Number0[23][5] = 4'hF;
    Number0[0][6] = 4'hF;
    Number0[1][6] = 4'hF;
    Number0[2][6] = 4'hF;
    Number0[3][6] = 4'hF;
    Number0[4][6] = 4'hF;
    Number0[5][6] = 4'hF;
    Number0[6][6] = 4'hF;
    Number0[7][6] = 4'hC;
    Number0[8][6] = 4'hC;
    Number0[9][6] = 4'hC;
    Number0[10][6] = 4'hC;
    Number0[11][6] = 4'hC;
    Number0[12][6] = 4'hC;
    Number0[13][6] = 4'hC;
    Number0[14][6] = 4'hC;
    Number0[15][6] = 4'hC;
    Number0[16][6] = 4'hC;
    Number0[17][6] = 4'hF;
    Number0[18][6] = 4'hF;
    Number0[19][6] = 4'hF;
    Number0[20][6] = 4'hF;
    Number0[21][6] = 4'hF;
    Number0[22][6] = 4'hF;
    Number0[23][6] = 4'hF;
    Number0[0][7] = 4'hF;
    Number0[1][7] = 4'hF;
    Number0[2][7] = 4'hF;
    Number0[3][7] = 4'hF;
    Number0[4][7] = 4'hF;
    Number0[5][7] = 4'hF;
    Number0[6][7] = 4'hF;
    Number0[7][7] = 4'hC;
    Number0[8][7] = 4'hC;
    Number0[9][7] = 4'hC;
    Number0[10][7] = 4'hC;
    Number0[11][7] = 4'hC;
    Number0[12][7] = 4'hC;
    Number0[13][7] = 4'hC;
    Number0[14][7] = 4'hC;
    Number0[15][7] = 4'hC;
    Number0[16][7] = 4'hC;
    Number0[17][7] = 4'hF;
    Number0[18][7] = 4'hF;
    Number0[19][7] = 4'hF;
    Number0[20][7] = 4'hF;
    Number0[21][7] = 4'hF;
    Number0[22][7] = 4'hF;
    Number0[23][7] = 4'hF;
    Number0[0][8] = 4'hF;
    Number0[1][8] = 4'hF;
    Number0[2][8] = 4'hC;
    Number0[3][8] = 4'hC;
    Number0[4][8] = 4'hC;
    Number0[5][8] = 4'hC;
    Number0[6][8] = 4'hC;
    Number0[7][8] = 4'hF;
    Number0[8][8] = 4'hF;
    Number0[9][8] = 4'hF;
    Number0[10][8] = 4'hF;
    Number0[11][8] = 4'hF;
    Number0[12][8] = 4'hF;
    Number0[13][8] = 4'hF;
    Number0[14][8] = 4'hF;
    Number0[15][8] = 4'hF;
    Number0[16][8] = 4'hF;
    Number0[17][8] = 4'hC;
    Number0[18][8] = 4'hC;
    Number0[19][8] = 4'hC;
    Number0[20][8] = 4'hC;
    Number0[21][8] = 4'hC;
    Number0[22][8] = 4'hF;
    Number0[23][8] = 4'hF;
    Number0[0][9] = 4'hF;
    Number0[1][9] = 4'hF;
    Number0[2][9] = 4'hC;
    Number0[3][9] = 4'hC;
    Number0[4][9] = 4'hC;
    Number0[5][9] = 4'hC;
    Number0[6][9] = 4'hC;
    Number0[7][9] = 4'hF;
    Number0[8][9] = 4'hF;
    Number0[9][9] = 4'hF;
    Number0[10][9] = 4'hF;
    Number0[11][9] = 4'hF;
    Number0[12][9] = 4'hF;
    Number0[13][9] = 4'hF;
    Number0[14][9] = 4'hF;
    Number0[15][9] = 4'hF;
    Number0[16][9] = 4'hF;
    Number0[17][9] = 4'hC;
    Number0[18][9] = 4'hC;
    Number0[19][9] = 4'hC;
    Number0[20][9] = 4'hC;
    Number0[21][9] = 4'hC;
    Number0[22][9] = 4'hF;
    Number0[23][9] = 4'hF;
    Number0[0][10] = 4'hF;
    Number0[1][10] = 4'hF;
    Number0[2][10] = 4'hC;
    Number0[3][10] = 4'hC;
    Number0[4][10] = 4'hC;
    Number0[5][10] = 4'hC;
    Number0[6][10] = 4'hC;
    Number0[7][10] = 4'hF;
    Number0[8][10] = 4'hF;
    Number0[9][10] = 4'hF;
    Number0[10][10] = 4'hF;
    Number0[11][10] = 4'hF;
    Number0[12][10] = 4'hF;
    Number0[13][10] = 4'hF;
    Number0[14][10] = 4'hF;
    Number0[15][10] = 4'hF;
    Number0[16][10] = 4'hF;
    Number0[17][10] = 4'hC;
    Number0[18][10] = 4'hC;
    Number0[19][10] = 4'hC;
    Number0[20][10] = 4'hC;
    Number0[21][10] = 4'hC;
    Number0[22][10] = 4'hF;
    Number0[23][10] = 4'hF;
    Number0[0][11] = 4'hF;
    Number0[1][11] = 4'hF;
    Number0[2][11] = 4'hC;
    Number0[3][11] = 4'hC;
    Number0[4][11] = 4'hC;
    Number0[5][11] = 4'hC;
    Number0[6][11] = 4'hC;
    Number0[7][11] = 4'hF;
    Number0[8][11] = 4'hF;
    Number0[9][11] = 4'hF;
    Number0[10][11] = 4'hF;
    Number0[11][11] = 4'hF;
    Number0[12][11] = 4'hF;
    Number0[13][11] = 4'hF;
    Number0[14][11] = 4'hF;
    Number0[15][11] = 4'hF;
    Number0[16][11] = 4'hF;
    Number0[17][11] = 4'hC;
    Number0[18][11] = 4'hC;
    Number0[19][11] = 4'hC;
    Number0[20][11] = 4'hC;
    Number0[21][11] = 4'hC;
    Number0[22][11] = 4'hF;
    Number0[23][11] = 4'hF;
    Number0[0][12] = 4'hF;
    Number0[1][12] = 4'hF;
    Number0[2][12] = 4'hC;
    Number0[3][12] = 4'hC;
    Number0[4][12] = 4'hC;
    Number0[5][12] = 4'hC;
    Number0[6][12] = 4'hC;
    Number0[7][12] = 4'hF;
    Number0[8][12] = 4'hF;
    Number0[9][12] = 4'hF;
    Number0[10][12] = 4'hF;
    Number0[11][12] = 4'hF;
    Number0[12][12] = 4'hF;
    Number0[13][12] = 4'hF;
    Number0[14][12] = 4'hF;
    Number0[15][12] = 4'hF;
    Number0[16][12] = 4'hF;
    Number0[17][12] = 4'hC;
    Number0[18][12] = 4'hC;
    Number0[19][12] = 4'hC;
    Number0[20][12] = 4'hC;
    Number0[21][12] = 4'hC;
    Number0[22][12] = 4'hF;
    Number0[23][12] = 4'hF;
    Number0[0][13] = 4'hF;
    Number0[1][13] = 4'hF;
    Number0[2][13] = 4'hC;
    Number0[3][13] = 4'hC;
    Number0[4][13] = 4'hC;
    Number0[5][13] = 4'hC;
    Number0[6][13] = 4'hC;
    Number0[7][13] = 4'hF;
    Number0[8][13] = 4'hF;
    Number0[9][13] = 4'hF;
    Number0[10][13] = 4'hF;
    Number0[11][13] = 4'hF;
    Number0[12][13] = 4'hF;
    Number0[13][13] = 4'hF;
    Number0[14][13] = 4'hF;
    Number0[15][13] = 4'hF;
    Number0[16][13] = 4'hF;
    Number0[17][13] = 4'hC;
    Number0[18][13] = 4'hC;
    Number0[19][13] = 4'hC;
    Number0[20][13] = 4'hC;
    Number0[21][13] = 4'hC;
    Number0[22][13] = 4'hF;
    Number0[23][13] = 4'hF;
    Number0[0][14] = 4'hF;
    Number0[1][14] = 4'hF;
    Number0[2][14] = 4'hC;
    Number0[3][14] = 4'hC;
    Number0[4][14] = 4'hC;
    Number0[5][14] = 4'hC;
    Number0[6][14] = 4'hC;
    Number0[7][14] = 4'hF;
    Number0[8][14] = 4'hF;
    Number0[9][14] = 4'hF;
    Number0[10][14] = 4'hF;
    Number0[11][14] = 4'hF;
    Number0[12][14] = 4'hF;
    Number0[13][14] = 4'hF;
    Number0[14][14] = 4'hF;
    Number0[15][14] = 4'hF;
    Number0[16][14] = 4'hF;
    Number0[17][14] = 4'hC;
    Number0[18][14] = 4'hC;
    Number0[19][14] = 4'hC;
    Number0[20][14] = 4'hC;
    Number0[21][14] = 4'hC;
    Number0[22][14] = 4'hF;
    Number0[23][14] = 4'hF;
    Number0[0][15] = 4'hF;
    Number0[1][15] = 4'hF;
    Number0[2][15] = 4'hC;
    Number0[3][15] = 4'hC;
    Number0[4][15] = 4'hC;
    Number0[5][15] = 4'hC;
    Number0[6][15] = 4'hC;
    Number0[7][15] = 4'hF;
    Number0[8][15] = 4'hF;
    Number0[9][15] = 4'hF;
    Number0[10][15] = 4'hF;
    Number0[11][15] = 4'hF;
    Number0[12][15] = 4'hF;
    Number0[13][15] = 4'hF;
    Number0[14][15] = 4'hF;
    Number0[15][15] = 4'hF;
    Number0[16][15] = 4'hF;
    Number0[17][15] = 4'hC;
    Number0[18][15] = 4'hC;
    Number0[19][15] = 4'hC;
    Number0[20][15] = 4'hC;
    Number0[21][15] = 4'hC;
    Number0[22][15] = 4'hF;
    Number0[23][15] = 4'hF;
    Number0[0][16] = 4'hF;
    Number0[1][16] = 4'hF;
    Number0[2][16] = 4'hC;
    Number0[3][16] = 4'hC;
    Number0[4][16] = 4'hC;
    Number0[5][16] = 4'hC;
    Number0[6][16] = 4'hC;
    Number0[7][16] = 4'hF;
    Number0[8][16] = 4'hF;
    Number0[9][16] = 4'hF;
    Number0[10][16] = 4'hF;
    Number0[11][16] = 4'hF;
    Number0[12][16] = 4'hF;
    Number0[13][16] = 4'hF;
    Number0[14][16] = 4'hF;
    Number0[15][16] = 4'hF;
    Number0[16][16] = 4'hF;
    Number0[17][16] = 4'hC;
    Number0[18][16] = 4'hC;
    Number0[19][16] = 4'hC;
    Number0[20][16] = 4'hC;
    Number0[21][16] = 4'hC;
    Number0[22][16] = 4'hF;
    Number0[23][16] = 4'hF;
    Number0[0][17] = 4'hF;
    Number0[1][17] = 4'hF;
    Number0[2][17] = 4'hC;
    Number0[3][17] = 4'hC;
    Number0[4][17] = 4'hC;
    Number0[5][17] = 4'hC;
    Number0[6][17] = 4'hC;
    Number0[7][17] = 4'hF;
    Number0[8][17] = 4'hF;
    Number0[9][17] = 4'hF;
    Number0[10][17] = 4'hF;
    Number0[11][17] = 4'hF;
    Number0[12][17] = 4'hF;
    Number0[13][17] = 4'hF;
    Number0[14][17] = 4'hF;
    Number0[15][17] = 4'hF;
    Number0[16][17] = 4'hF;
    Number0[17][17] = 4'hC;
    Number0[18][17] = 4'hC;
    Number0[19][17] = 4'hC;
    Number0[20][17] = 4'hC;
    Number0[21][17] = 4'hC;
    Number0[22][17] = 4'hF;
    Number0[23][17] = 4'hF;
    Number0[0][18] = 4'hF;
    Number0[1][18] = 4'hF;
    Number0[2][18] = 4'hC;
    Number0[3][18] = 4'hC;
    Number0[4][18] = 4'hC;
    Number0[5][18] = 4'hC;
    Number0[6][18] = 4'hC;
    Number0[7][18] = 4'hF;
    Number0[8][18] = 4'hF;
    Number0[9][18] = 4'hF;
    Number0[10][18] = 4'hF;
    Number0[11][18] = 4'hF;
    Number0[12][18] = 4'hF;
    Number0[13][18] = 4'hF;
    Number0[14][18] = 4'hF;
    Number0[15][18] = 4'hF;
    Number0[16][18] = 4'hF;
    Number0[17][18] = 4'hC;
    Number0[18][18] = 4'hC;
    Number0[19][18] = 4'hC;
    Number0[20][18] = 4'hC;
    Number0[21][18] = 4'hC;
    Number0[22][18] = 4'hF;
    Number0[23][18] = 4'hF;
    Number0[0][19] = 4'hF;
    Number0[1][19] = 4'hF;
    Number0[2][19] = 4'hC;
    Number0[3][19] = 4'hC;
    Number0[4][19] = 4'hC;
    Number0[5][19] = 4'hC;
    Number0[6][19] = 4'hC;
    Number0[7][19] = 4'hF;
    Number0[8][19] = 4'hF;
    Number0[9][19] = 4'hF;
    Number0[10][19] = 4'hF;
    Number0[11][19] = 4'hF;
    Number0[12][19] = 4'hF;
    Number0[13][19] = 4'hF;
    Number0[14][19] = 4'hF;
    Number0[15][19] = 4'hF;
    Number0[16][19] = 4'hF;
    Number0[17][19] = 4'hC;
    Number0[18][19] = 4'hC;
    Number0[19][19] = 4'hC;
    Number0[20][19] = 4'hC;
    Number0[21][19] = 4'hC;
    Number0[22][19] = 4'hF;
    Number0[23][19] = 4'hF;
    Number0[0][20] = 4'hF;
    Number0[1][20] = 4'hF;
    Number0[2][20] = 4'hC;
    Number0[3][20] = 4'hC;
    Number0[4][20] = 4'hC;
    Number0[5][20] = 4'hC;
    Number0[6][20] = 4'hC;
    Number0[7][20] = 4'hF;
    Number0[8][20] = 4'hF;
    Number0[9][20] = 4'hF;
    Number0[10][20] = 4'hF;
    Number0[11][20] = 4'hF;
    Number0[12][20] = 4'hF;
    Number0[13][20] = 4'hF;
    Number0[14][20] = 4'hF;
    Number0[15][20] = 4'hF;
    Number0[16][20] = 4'hF;
    Number0[17][20] = 4'hC;
    Number0[18][20] = 4'hC;
    Number0[19][20] = 4'hC;
    Number0[20][20] = 4'hC;
    Number0[21][20] = 4'hC;
    Number0[22][20] = 4'hF;
    Number0[23][20] = 4'hF;
    Number0[0][21] = 4'hF;
    Number0[1][21] = 4'hF;
    Number0[2][21] = 4'hC;
    Number0[3][21] = 4'hC;
    Number0[4][21] = 4'hC;
    Number0[5][21] = 4'hC;
    Number0[6][21] = 4'hC;
    Number0[7][21] = 4'hF;
    Number0[8][21] = 4'hF;
    Number0[9][21] = 4'hF;
    Number0[10][21] = 4'hF;
    Number0[11][21] = 4'hF;
    Number0[12][21] = 4'hF;
    Number0[13][21] = 4'hF;
    Number0[14][21] = 4'hF;
    Number0[15][21] = 4'hF;
    Number0[16][21] = 4'hF;
    Number0[17][21] = 4'hC;
    Number0[18][21] = 4'hC;
    Number0[19][21] = 4'hC;
    Number0[20][21] = 4'hC;
    Number0[21][21] = 4'hC;
    Number0[22][21] = 4'hF;
    Number0[23][21] = 4'hF;
    Number0[0][22] = 4'hF;
    Number0[1][22] = 4'hF;
    Number0[2][22] = 4'hC;
    Number0[3][22] = 4'hC;
    Number0[4][22] = 4'hC;
    Number0[5][22] = 4'hC;
    Number0[6][22] = 4'hC;
    Number0[7][22] = 4'hF;
    Number0[8][22] = 4'hF;
    Number0[9][22] = 4'hF;
    Number0[10][22] = 4'hF;
    Number0[11][22] = 4'hF;
    Number0[12][22] = 4'hF;
    Number0[13][22] = 4'hF;
    Number0[14][22] = 4'hF;
    Number0[15][22] = 4'hF;
    Number0[16][22] = 4'hF;
    Number0[17][22] = 4'hC;
    Number0[18][22] = 4'hC;
    Number0[19][22] = 4'hC;
    Number0[20][22] = 4'hC;
    Number0[21][22] = 4'hC;
    Number0[22][22] = 4'hF;
    Number0[23][22] = 4'hF;
    Number0[0][23] = 4'hF;
    Number0[1][23] = 4'hF;
    Number0[2][23] = 4'hF;
    Number0[3][23] = 4'hF;
    Number0[4][23] = 4'hF;
    Number0[5][23] = 4'hF;
    Number0[6][23] = 4'hF;
    Number0[7][23] = 4'hC;
    Number0[8][23] = 4'hC;
    Number0[9][23] = 4'hC;
    Number0[10][23] = 4'hC;
    Number0[11][23] = 4'hC;
    Number0[12][23] = 4'hC;
    Number0[13][23] = 4'hC;
    Number0[14][23] = 4'hC;
    Number0[15][23] = 4'hC;
    Number0[16][23] = 4'hC;
    Number0[17][23] = 4'hF;
    Number0[18][23] = 4'hF;
    Number0[19][23] = 4'hF;
    Number0[20][23] = 4'hF;
    Number0[21][23] = 4'hF;
    Number0[22][23] = 4'hF;
    Number0[23][23] = 4'hF;
    Number0[0][24] = 4'hF;
    Number0[1][24] = 4'hF;
    Number0[2][24] = 4'hF;
    Number0[3][24] = 4'hF;
    Number0[4][24] = 4'hF;
    Number0[5][24] = 4'hF;
    Number0[6][24] = 4'hF;
    Number0[7][24] = 4'hC;
    Number0[8][24] = 4'hC;
    Number0[9][24] = 4'hC;
    Number0[10][24] = 4'hC;
    Number0[11][24] = 4'hC;
    Number0[12][24] = 4'hC;
    Number0[13][24] = 4'hC;
    Number0[14][24] = 4'hC;
    Number0[15][24] = 4'hC;
    Number0[16][24] = 4'hC;
    Number0[17][24] = 4'hF;
    Number0[18][24] = 4'hF;
    Number0[19][24] = 4'hF;
    Number0[20][24] = 4'hF;
    Number0[21][24] = 4'hF;
    Number0[22][24] = 4'hF;
    Number0[23][24] = 4'hF;
    Number0[0][25] = 4'hF;
    Number0[1][25] = 4'hF;
    Number0[2][25] = 4'hF;
    Number0[3][25] = 4'hF;
    Number0[4][25] = 4'hF;
    Number0[5][25] = 4'hF;
    Number0[6][25] = 4'hF;
    Number0[7][25] = 4'hC;
    Number0[8][25] = 4'hC;
    Number0[9][25] = 4'hC;
    Number0[10][25] = 4'hC;
    Number0[11][25] = 4'hC;
    Number0[12][25] = 4'hC;
    Number0[13][25] = 4'hC;
    Number0[14][25] = 4'hC;
    Number0[15][25] = 4'hC;
    Number0[16][25] = 4'hC;
    Number0[17][25] = 4'hF;
    Number0[18][25] = 4'hF;
    Number0[19][25] = 4'hF;
    Number0[20][25] = 4'hF;
    Number0[21][25] = 4'hF;
    Number0[22][25] = 4'hF;
    Number0[23][25] = 4'hF;
    Number0[0][26] = 4'hF;
    Number0[1][26] = 4'hF;
    Number0[2][26] = 4'hF;
    Number0[3][26] = 4'hF;
    Number0[4][26] = 4'hF;
    Number0[5][26] = 4'hF;
    Number0[6][26] = 4'hF;
    Number0[7][26] = 4'hC;
    Number0[8][26] = 4'hC;
    Number0[9][26] = 4'hC;
    Number0[10][26] = 4'hC;
    Number0[11][26] = 4'hC;
    Number0[12][26] = 4'hC;
    Number0[13][26] = 4'hC;
    Number0[14][26] = 4'hC;
    Number0[15][26] = 4'hC;
    Number0[16][26] = 4'hC;
    Number0[17][26] = 4'hF;
    Number0[18][26] = 4'hF;
    Number0[19][26] = 4'hF;
    Number0[20][26] = 4'hF;
    Number0[21][26] = 4'hF;
    Number0[22][26] = 4'hF;
    Number0[23][26] = 4'hF;
    Number0[0][27] = 4'hF;
    Number0[1][27] = 4'hF;
    Number0[2][27] = 4'hF;
    Number0[3][27] = 4'hF;
    Number0[4][27] = 4'hF;
    Number0[5][27] = 4'hF;
    Number0[6][27] = 4'hF;
    Number0[7][27] = 4'hC;
    Number0[8][27] = 4'hC;
    Number0[9][27] = 4'hC;
    Number0[10][27] = 4'hC;
    Number0[11][27] = 4'hC;
    Number0[12][27] = 4'hC;
    Number0[13][27] = 4'hC;
    Number0[14][27] = 4'hC;
    Number0[15][27] = 4'hC;
    Number0[16][27] = 4'hC;
    Number0[17][27] = 4'hF;
    Number0[18][27] = 4'hF;
    Number0[19][27] = 4'hF;
    Number0[20][27] = 4'hF;
    Number0[21][27] = 4'hF;
    Number0[22][27] = 4'hF;
    Number0[23][27] = 4'hF;
    Number0[0][28] = 4'hF;
    Number0[1][28] = 4'hF;
    Number0[2][28] = 4'hF;
    Number0[3][28] = 4'hF;
    Number0[4][28] = 4'hF;
    Number0[5][28] = 4'hF;
    Number0[6][28] = 4'hF;
    Number0[7][28] = 4'hF;
    Number0[8][28] = 4'hF;
    Number0[9][28] = 4'hF;
    Number0[10][28] = 4'hF;
    Number0[11][28] = 4'hF;
    Number0[12][28] = 4'hF;
    Number0[13][28] = 4'hF;
    Number0[14][28] = 4'hF;
    Number0[15][28] = 4'hF;
    Number0[16][28] = 4'hF;
    Number0[17][28] = 4'hF;
    Number0[18][28] = 4'hF;
    Number0[19][28] = 4'hF;
    Number0[20][28] = 4'hF;
    Number0[21][28] = 4'hF;
    Number0[22][28] = 4'hF;
    Number0[23][28] = 4'hF;
    Number0[0][29] = 4'hF;
    Number0[1][29] = 4'hF;
    Number0[2][29] = 4'hF;
    Number0[3][29] = 4'hF;
    Number0[4][29] = 4'hF;
    Number0[5][29] = 4'hF;
    Number0[6][29] = 4'hF;
    Number0[7][29] = 4'hF;
    Number0[8][29] = 4'hF;
    Number0[9][29] = 4'hF;
    Number0[10][29] = 4'hF;
    Number0[11][29] = 4'hF;
    Number0[12][29] = 4'hF;
    Number0[13][29] = 4'hF;
    Number0[14][29] = 4'hF;
    Number0[15][29] = 4'hF;
    Number0[16][29] = 4'hF;
    Number0[17][29] = 4'hF;
    Number0[18][29] = 4'hF;
    Number0[19][29] = 4'hF;
    Number0[20][29] = 4'hF;
    Number0[21][29] = 4'hF;
    Number0[22][29] = 4'hF;
    Number0[23][29] = 4'hF;
 
//Number 1
    Number1[0][0] = 4'hF;
    Number1[1][0] = 4'hF;
    Number1[2][0] = 4'hF;
    Number1[3][0] = 4'hF;
    Number1[4][0] = 4'hF;
    Number1[5][0] = 4'hF;
    Number1[6][0] = 4'hF;
    Number1[7][0] = 4'hF;
    Number1[8][0] = 4'hF;
    Number1[9][0] = 4'hF;
    Number1[10][0] = 4'hF;
    Number1[11][0] = 4'hF;
    Number1[12][0] = 4'hF;
    Number1[13][0] = 4'hF;
    Number1[14][0] = 4'hF;
    Number1[15][0] = 4'hF;
    Number1[16][0] = 4'hF;
    Number1[17][0] = 4'hF;
    Number1[18][0] = 4'hF;
    Number1[19][0] = 4'hF;
    Number1[20][0] = 4'hF;
    Number1[21][0] = 4'hF;
    Number1[22][0] = 4'hF;
    Number1[23][0] = 4'hF;
    Number1[0][1] = 4'hF;
    Number1[1][1] = 4'hF;
    Number1[2][1] = 4'hF;
    Number1[3][1] = 4'hF;
    Number1[4][1] = 4'hF;
    Number1[5][1] = 4'hF;
    Number1[6][1] = 4'hF;
    Number1[7][1] = 4'hF;
    Number1[8][1] = 4'hF;
    Number1[9][1] = 4'hF;
    Number1[10][1] = 4'hF;
    Number1[11][1] = 4'hF;
    Number1[12][1] = 4'hF;
    Number1[13][1] = 4'hF;
    Number1[14][1] = 4'hF;
    Number1[15][1] = 4'hF;
    Number1[16][1] = 4'hF;
    Number1[17][1] = 4'hF;
    Number1[18][1] = 4'hF;
    Number1[19][1] = 4'hF;
    Number1[20][1] = 4'hF;
    Number1[21][1] = 4'hF;
    Number1[22][1] = 4'hF;
    Number1[23][1] = 4'hF;
    Number1[0][2] = 4'hF;
    Number1[1][2] = 4'hF;
    Number1[2][2] = 4'hF;
    Number1[3][2] = 4'hF;
    Number1[4][2] = 4'hF;
    Number1[5][2] = 4'hF;
    Number1[6][2] = 4'hF;
    Number1[7][2] = 4'hF;
    Number1[8][2] = 4'hF;
    Number1[9][2] = 4'hF;
    Number1[10][2] = 4'hF;
    Number1[11][2] = 4'hF;
    Number1[12][2] = 4'hF;
    Number1[13][2] = 4'hF;
    Number1[14][2] = 4'hF;
    Number1[15][2] = 4'hF;
    Number1[16][2] = 4'hF;
    Number1[17][2] = 4'hF;
    Number1[18][2] = 4'hF;
    Number1[19][2] = 4'hF;
    Number1[20][2] = 4'hF;
    Number1[21][2] = 4'hF;
    Number1[22][2] = 4'hF;
    Number1[23][2] = 4'hF;
    Number1[0][3] = 4'hF;
    Number1[1][3] = 4'hF;
    Number1[2][3] = 4'hF;
    Number1[3][3] = 4'hF;
    Number1[4][3] = 4'hF;
    Number1[5][3] = 4'hF;
    Number1[6][3] = 4'hF;
    Number1[7][3] = 4'hC;
    Number1[8][3] = 4'hC;
    Number1[9][3] = 4'hC;
    Number1[10][3] = 4'hC;
    Number1[11][3] = 4'hC;
    Number1[12][3] = 4'hC;
    Number1[13][3] = 4'hC;
    Number1[14][3] = 4'hC;
    Number1[15][3] = 4'hC;
    Number1[16][3] = 4'hC;
    Number1[17][3] = 4'hF;
    Number1[18][3] = 4'hF;
    Number1[19][3] = 4'hF;
    Number1[20][3] = 4'hF;
    Number1[21][3] = 4'hF;
    Number1[22][3] = 4'hF;
    Number1[23][3] = 4'hF;
    Number1[0][4] = 4'hF;
    Number1[1][4] = 4'hF;
    Number1[2][4] = 4'hF;
    Number1[3][4] = 4'hF;
    Number1[4][4] = 4'hF;
    Number1[5][4] = 4'hF;
    Number1[6][4] = 4'hF;
    Number1[7][4] = 4'hC;
    Number1[8][4] = 4'hC;
    Number1[9][4] = 4'hC;
    Number1[10][4] = 4'hC;
    Number1[11][4] = 4'hC;
    Number1[12][4] = 4'hC;
    Number1[13][4] = 4'hC;
    Number1[14][4] = 4'hC;
    Number1[15][4] = 4'hC;
    Number1[16][4] = 4'hC;
    Number1[17][4] = 4'hF;
    Number1[18][4] = 4'hF;
    Number1[19][4] = 4'hF;
    Number1[20][4] = 4'hF;
    Number1[21][4] = 4'hF;
    Number1[22][4] = 4'hF;
    Number1[23][4] = 4'hF;
    Number1[0][5] = 4'hF;
    Number1[1][5] = 4'hF;
    Number1[2][5] = 4'hF;
    Number1[3][5] = 4'hF;
    Number1[4][5] = 4'hF;
    Number1[5][5] = 4'hF;
    Number1[6][5] = 4'hF;
    Number1[7][5] = 4'hC;
    Number1[8][5] = 4'hC;
    Number1[9][5] = 4'hC;
    Number1[10][5] = 4'hC;
    Number1[11][5] = 4'hC;
    Number1[12][5] = 4'hC;
    Number1[13][5] = 4'hC;
    Number1[14][5] = 4'hC;
    Number1[15][5] = 4'hC;
    Number1[16][5] = 4'hC;
    Number1[17][5] = 4'hF;
    Number1[18][5] = 4'hF;
    Number1[19][5] = 4'hF;
    Number1[20][5] = 4'hF;
    Number1[21][5] = 4'hF;
    Number1[22][5] = 4'hF;
    Number1[23][5] = 4'hF;
    Number1[0][6] = 4'hF;
    Number1[1][6] = 4'hF;
    Number1[2][6] = 4'hF;
    Number1[3][6] = 4'hF;
    Number1[4][6] = 4'hF;
    Number1[5][6] = 4'hF;
    Number1[6][6] = 4'hF;
    Number1[7][6] = 4'hC;
    Number1[8][6] = 4'hC;
    Number1[9][6] = 4'hC;
    Number1[10][6] = 4'hC;
    Number1[11][6] = 4'hC;
    Number1[12][6] = 4'hC;
    Number1[13][6] = 4'hC;
    Number1[14][6] = 4'hC;
    Number1[15][6] = 4'hC;
    Number1[16][6] = 4'hC;
    Number1[17][6] = 4'hF;
    Number1[18][6] = 4'hF;
    Number1[19][6] = 4'hF;
    Number1[20][6] = 4'hF;
    Number1[21][6] = 4'hF;
    Number1[22][6] = 4'hF;
    Number1[23][6] = 4'hF;
    Number1[0][7] = 4'hF;
    Number1[1][7] = 4'hF;
    Number1[2][7] = 4'hF;
    Number1[3][7] = 4'hF;
    Number1[4][7] = 4'hF;
    Number1[5][7] = 4'hF;
    Number1[6][7] = 4'hF;
    Number1[7][7] = 4'hC;
    Number1[8][7] = 4'hC;
    Number1[9][7] = 4'hC;
    Number1[10][7] = 4'hC;
    Number1[11][7] = 4'hC;
    Number1[12][7] = 4'hC;
    Number1[13][7] = 4'hC;
    Number1[14][7] = 4'hC;
    Number1[15][7] = 4'hC;
    Number1[16][7] = 4'hC;
    Number1[17][7] = 4'hF;
    Number1[18][7] = 4'hF;
    Number1[19][7] = 4'hF;
    Number1[20][7] = 4'hF;
    Number1[21][7] = 4'hF;
    Number1[22][7] = 4'hF;
    Number1[23][7] = 4'hF;
    Number1[0][8] = 4'hF;
    Number1[1][8] = 4'hF;
    Number1[2][8] = 4'hF;
    Number1[3][8] = 4'hF;
    Number1[4][8] = 4'hF;
    Number1[5][8] = 4'hF;
    Number1[6][8] = 4'hF;
    Number1[7][8] = 4'hF;
    Number1[8][8] = 4'hF;
    Number1[9][8] = 4'hF;
    Number1[10][8] = 4'hF;
    Number1[11][8] = 4'hF;
    Number1[12][8] = 4'hC;
    Number1[13][8] = 4'hC;
    Number1[14][8] = 4'hC;
    Number1[15][8] = 4'hC;
    Number1[16][8] = 4'hC;
    Number1[17][8] = 4'hF;
    Number1[18][8] = 4'hF;
    Number1[19][8] = 4'hF;
    Number1[20][8] = 4'hF;
    Number1[21][8] = 4'hF;
    Number1[22][8] = 4'hF;
    Number1[23][8] = 4'hF;
    Number1[0][9] = 4'hF;
    Number1[1][9] = 4'hF;
    Number1[2][9] = 4'hF;
    Number1[3][9] = 4'hF;
    Number1[4][9] = 4'hF;
    Number1[5][9] = 4'hF;
    Number1[6][9] = 4'hF;
    Number1[7][9] = 4'hF;
    Number1[8][9] = 4'hF;
    Number1[9][9] = 4'hF;
    Number1[10][9] = 4'hF;
    Number1[11][9] = 4'hF;
    Number1[12][9] = 4'hC;
    Number1[13][9] = 4'hC;
    Number1[14][9] = 4'hC;
    Number1[15][9] = 4'hC;
    Number1[16][9] = 4'hC;
    Number1[17][9] = 4'hF;
    Number1[18][9] = 4'hF;
    Number1[19][9] = 4'hF;
    Number1[20][9] = 4'hF;
    Number1[21][9] = 4'hF;
    Number1[22][9] = 4'hF;
    Number1[23][9] = 4'hF;
    Number1[0][10] = 4'hF;
    Number1[1][10] = 4'hF;
    Number1[2][10] = 4'hF;
    Number1[3][10] = 4'hF;
    Number1[4][10] = 4'hF;
    Number1[5][10] = 4'hF;
    Number1[6][10] = 4'hF;
    Number1[7][10] = 4'hF;
    Number1[8][10] = 4'hF;
    Number1[9][10] = 4'hF;
    Number1[10][10] = 4'hF;
    Number1[11][10] = 4'hF;
    Number1[12][10] = 4'hC;
    Number1[13][10] = 4'hC;
    Number1[14][10] = 4'hC;
    Number1[15][10] = 4'hC;
    Number1[16][10] = 4'hC;
    Number1[17][10] = 4'hF;
    Number1[18][10] = 4'hF;
    Number1[19][10] = 4'hF;
    Number1[20][10] = 4'hF;
    Number1[21][10] = 4'hF;
    Number1[22][10] = 4'hF;
    Number1[23][10] = 4'hF;
    Number1[0][11] = 4'hF;
    Number1[1][11] = 4'hF;
    Number1[2][11] = 4'hF;
    Number1[3][11] = 4'hF;
    Number1[4][11] = 4'hF;
    Number1[5][11] = 4'hF;
    Number1[6][11] = 4'hF;
    Number1[7][11] = 4'hF;
    Number1[8][11] = 4'hF;
    Number1[9][11] = 4'hF;
    Number1[10][11] = 4'hF;
    Number1[11][11] = 4'hF;
    Number1[12][11] = 4'hC;
    Number1[13][11] = 4'hC;
    Number1[14][11] = 4'hC;
    Number1[15][11] = 4'hC;
    Number1[16][11] = 4'hC;
    Number1[17][11] = 4'hF;
    Number1[18][11] = 4'hF;
    Number1[19][11] = 4'hF;
    Number1[20][11] = 4'hF;
    Number1[21][11] = 4'hF;
    Number1[22][11] = 4'hF;
    Number1[23][11] = 4'hF;
    Number1[0][12] = 4'hF;
    Number1[1][12] = 4'hF;
    Number1[2][12] = 4'hF;
    Number1[3][12] = 4'hF;
    Number1[4][12] = 4'hF;
    Number1[5][12] = 4'hF;
    Number1[6][12] = 4'hF;
    Number1[7][12] = 4'hF;
    Number1[8][12] = 4'hF;
    Number1[9][12] = 4'hF;
    Number1[10][12] = 4'hF;
    Number1[11][12] = 4'hF;
    Number1[12][12] = 4'hC;
    Number1[13][12] = 4'hC;
    Number1[14][12] = 4'hC;
    Number1[15][12] = 4'hC;
    Number1[16][12] = 4'hC;
    Number1[17][12] = 4'hF;
    Number1[18][12] = 4'hF;
    Number1[19][12] = 4'hF;
    Number1[20][12] = 4'hF;
    Number1[21][12] = 4'hF;
    Number1[22][12] = 4'hF;
    Number1[23][12] = 4'hF;
    Number1[0][13] = 4'hF;
    Number1[1][13] = 4'hF;
    Number1[2][13] = 4'hF;
    Number1[3][13] = 4'hF;
    Number1[4][13] = 4'hF;
    Number1[5][13] = 4'hF;
    Number1[6][13] = 4'hF;
    Number1[7][13] = 4'hF;
    Number1[8][13] = 4'hF;
    Number1[9][13] = 4'hF;
    Number1[10][13] = 4'hF;
    Number1[11][13] = 4'hF;
    Number1[12][13] = 4'hC;
    Number1[13][13] = 4'hC;
    Number1[14][13] = 4'hC;
    Number1[15][13] = 4'hC;
    Number1[16][13] = 4'hC;
    Number1[17][13] = 4'hF;
    Number1[18][13] = 4'hF;
    Number1[19][13] = 4'hF;
    Number1[20][13] = 4'hF;
    Number1[21][13] = 4'hF;
    Number1[22][13] = 4'hF;
    Number1[23][13] = 4'hF;
    Number1[0][14] = 4'hF;
    Number1[1][14] = 4'hF;
    Number1[2][14] = 4'hF;
    Number1[3][14] = 4'hF;
    Number1[4][14] = 4'hF;
    Number1[5][14] = 4'hF;
    Number1[6][14] = 4'hF;
    Number1[7][14] = 4'hF;
    Number1[8][14] = 4'hF;
    Number1[9][14] = 4'hF;
    Number1[10][14] = 4'hF;
    Number1[11][14] = 4'hF;
    Number1[12][14] = 4'hC;
    Number1[13][14] = 4'hC;
    Number1[14][14] = 4'hC;
    Number1[15][14] = 4'hC;
    Number1[16][14] = 4'hC;
    Number1[17][14] = 4'hF;
    Number1[18][14] = 4'hF;
    Number1[19][14] = 4'hF;
    Number1[20][14] = 4'hF;
    Number1[21][14] = 4'hF;
    Number1[22][14] = 4'hF;
    Number1[23][14] = 4'hF;
    Number1[0][15] = 4'hF;
    Number1[1][15] = 4'hF;
    Number1[2][15] = 4'hF;
    Number1[3][15] = 4'hF;
    Number1[4][15] = 4'hF;
    Number1[5][15] = 4'hF;
    Number1[6][15] = 4'hF;
    Number1[7][15] = 4'hF;
    Number1[8][15] = 4'hF;
    Number1[9][15] = 4'hF;
    Number1[10][15] = 4'hF;
    Number1[11][15] = 4'hF;
    Number1[12][15] = 4'hC;
    Number1[13][15] = 4'hC;
    Number1[14][15] = 4'hC;
    Number1[15][15] = 4'hC;
    Number1[16][15] = 4'hC;
    Number1[17][15] = 4'hF;
    Number1[18][15] = 4'hF;
    Number1[19][15] = 4'hF;
    Number1[20][15] = 4'hF;
    Number1[21][15] = 4'hF;
    Number1[22][15] = 4'hF;
    Number1[23][15] = 4'hF;
    Number1[0][16] = 4'hF;
    Number1[1][16] = 4'hF;
    Number1[2][16] = 4'hF;
    Number1[3][16] = 4'hF;
    Number1[4][16] = 4'hF;
    Number1[5][16] = 4'hF;
    Number1[6][16] = 4'hF;
    Number1[7][16] = 4'hF;
    Number1[8][16] = 4'hF;
    Number1[9][16] = 4'hF;
    Number1[10][16] = 4'hF;
    Number1[11][16] = 4'hF;
    Number1[12][16] = 4'hC;
    Number1[13][16] = 4'hC;
    Number1[14][16] = 4'hC;
    Number1[15][16] = 4'hC;
    Number1[16][16] = 4'hC;
    Number1[17][16] = 4'hF;
    Number1[18][16] = 4'hF;
    Number1[19][16] = 4'hF;
    Number1[20][16] = 4'hF;
    Number1[21][16] = 4'hF;
    Number1[22][16] = 4'hF;
    Number1[23][16] = 4'hF;
    Number1[0][17] = 4'hF;
    Number1[1][17] = 4'hF;
    Number1[2][17] = 4'hF;
    Number1[3][17] = 4'hF;
    Number1[4][17] = 4'hF;
    Number1[5][17] = 4'hF;
    Number1[6][17] = 4'hF;
    Number1[7][17] = 4'hF;
    Number1[8][17] = 4'hF;
    Number1[9][17] = 4'hF;
    Number1[10][17] = 4'hF;
    Number1[11][17] = 4'hF;
    Number1[12][17] = 4'hC;
    Number1[13][17] = 4'hC;
    Number1[14][17] = 4'hC;
    Number1[15][17] = 4'hC;
    Number1[16][17] = 4'hC;
    Number1[17][17] = 4'hF;
    Number1[18][17] = 4'hF;
    Number1[19][17] = 4'hF;
    Number1[20][17] = 4'hF;
    Number1[21][17] = 4'hF;
    Number1[22][17] = 4'hF;
    Number1[23][17] = 4'hF;
    Number1[0][18] = 4'hF;
    Number1[1][18] = 4'hF;
    Number1[2][18] = 4'hF;
    Number1[3][18] = 4'hF;
    Number1[4][18] = 4'hF;
    Number1[5][18] = 4'hF;
    Number1[6][18] = 4'hF;
    Number1[7][18] = 4'hF;
    Number1[8][18] = 4'hF;
    Number1[9][18] = 4'hF;
    Number1[10][18] = 4'hF;
    Number1[11][18] = 4'hF;
    Number1[12][18] = 4'hC;
    Number1[13][18] = 4'hC;
    Number1[14][18] = 4'hC;
    Number1[15][18] = 4'hC;
    Number1[16][18] = 4'hC;
    Number1[17][18] = 4'hF;
    Number1[18][18] = 4'hF;
    Number1[19][18] = 4'hF;
    Number1[20][18] = 4'hF;
    Number1[21][18] = 4'hF;
    Number1[22][18] = 4'hF;
    Number1[23][18] = 4'hF;
    Number1[0][19] = 4'hF;
    Number1[1][19] = 4'hF;
    Number1[2][19] = 4'hF;
    Number1[3][19] = 4'hF;
    Number1[4][19] = 4'hF;
    Number1[5][19] = 4'hF;
    Number1[6][19] = 4'hF;
    Number1[7][19] = 4'hF;
    Number1[8][19] = 4'hF;
    Number1[9][19] = 4'hF;
    Number1[10][19] = 4'hF;
    Number1[11][19] = 4'hF;
    Number1[12][19] = 4'hC;
    Number1[13][19] = 4'hC;
    Number1[14][19] = 4'hC;
    Number1[15][19] = 4'hC;
    Number1[16][19] = 4'hC;
    Number1[17][19] = 4'hF;
    Number1[18][19] = 4'hF;
    Number1[19][19] = 4'hF;
    Number1[20][19] = 4'hF;
    Number1[21][19] = 4'hF;
    Number1[22][19] = 4'hF;
    Number1[23][19] = 4'hF;
    Number1[0][20] = 4'hF;
    Number1[1][20] = 4'hF;
    Number1[2][20] = 4'hF;
    Number1[3][20] = 4'hF;
    Number1[4][20] = 4'hF;
    Number1[5][20] = 4'hF;
    Number1[6][20] = 4'hF;
    Number1[7][20] = 4'hF;
    Number1[8][20] = 4'hF;
    Number1[9][20] = 4'hF;
    Number1[10][20] = 4'hF;
    Number1[11][20] = 4'hF;
    Number1[12][20] = 4'hC;
    Number1[13][20] = 4'hC;
    Number1[14][20] = 4'hC;
    Number1[15][20] = 4'hC;
    Number1[16][20] = 4'hC;
    Number1[17][20] = 4'hF;
    Number1[18][20] = 4'hF;
    Number1[19][20] = 4'hF;
    Number1[20][20] = 4'hF;
    Number1[21][20] = 4'hF;
    Number1[22][20] = 4'hF;
    Number1[23][20] = 4'hF;
    Number1[0][21] = 4'hF;
    Number1[1][21] = 4'hF;
    Number1[2][21] = 4'hF;
    Number1[3][21] = 4'hF;
    Number1[4][21] = 4'hF;
    Number1[5][21] = 4'hF;
    Number1[6][21] = 4'hF;
    Number1[7][21] = 4'hF;
    Number1[8][21] = 4'hF;
    Number1[9][21] = 4'hF;
    Number1[10][21] = 4'hF;
    Number1[11][21] = 4'hF;
    Number1[12][21] = 4'hC;
    Number1[13][21] = 4'hC;
    Number1[14][21] = 4'hC;
    Number1[15][21] = 4'hC;
    Number1[16][21] = 4'hC;
    Number1[17][21] = 4'hF;
    Number1[18][21] = 4'hF;
    Number1[19][21] = 4'hF;
    Number1[20][21] = 4'hF;
    Number1[21][21] = 4'hF;
    Number1[22][21] = 4'hF;
    Number1[23][21] = 4'hF;
    Number1[0][22] = 4'hF;
    Number1[1][22] = 4'hF;
    Number1[2][22] = 4'hF;
    Number1[3][22] = 4'hF;
    Number1[4][22] = 4'hF;
    Number1[5][22] = 4'hF;
    Number1[6][22] = 4'hF;
    Number1[7][22] = 4'hF;
    Number1[8][22] = 4'hF;
    Number1[9][22] = 4'hF;
    Number1[10][22] = 4'hF;
    Number1[11][22] = 4'hF;
    Number1[12][22] = 4'hC;
    Number1[13][22] = 4'hC;
    Number1[14][22] = 4'hC;
    Number1[15][22] = 4'hC;
    Number1[16][22] = 4'hC;
    Number1[17][22] = 4'hF;
    Number1[18][22] = 4'hF;
    Number1[19][22] = 4'hF;
    Number1[20][22] = 4'hF;
    Number1[21][22] = 4'hF;
    Number1[22][22] = 4'hF;
    Number1[23][22] = 4'hF;
    Number1[0][23] = 4'hF;
    Number1[1][23] = 4'hF;
    Number1[2][23] = 4'hF;
    Number1[3][23] = 4'hF;
    Number1[4][23] = 4'hF;
    Number1[5][23] = 4'hF;
    Number1[6][23] = 4'hF;
    Number1[7][23] = 4'hF;
    Number1[8][23] = 4'hF;
    Number1[9][23] = 4'hF;
    Number1[10][23] = 4'hF;
    Number1[11][23] = 4'hF;
    Number1[12][23] = 4'hC;
    Number1[13][23] = 4'hC;
    Number1[14][23] = 4'hC;
    Number1[15][23] = 4'hC;
    Number1[16][23] = 4'hC;
    Number1[17][23] = 4'hF;
    Number1[18][23] = 4'hF;
    Number1[19][23] = 4'hF;
    Number1[20][23] = 4'hF;
    Number1[21][23] = 4'hF;
    Number1[22][23] = 4'hF;
    Number1[23][23] = 4'hF;
    Number1[0][24] = 4'hF;
    Number1[1][24] = 4'hF;
    Number1[2][24] = 4'hF;
    Number1[3][24] = 4'hF;
    Number1[4][24] = 4'hF;
    Number1[5][24] = 4'hF;
    Number1[6][24] = 4'hF;
    Number1[7][24] = 4'hF;
    Number1[8][24] = 4'hF;
    Number1[9][24] = 4'hF;
    Number1[10][24] = 4'hF;
    Number1[11][24] = 4'hF;
    Number1[12][24] = 4'hC;
    Number1[13][24] = 4'hC;
    Number1[14][24] = 4'hC;
    Number1[15][24] = 4'hC;
    Number1[16][24] = 4'hC;
    Number1[17][24] = 4'hF;
    Number1[18][24] = 4'hF;
    Number1[19][24] = 4'hF;
    Number1[20][24] = 4'hF;
    Number1[21][24] = 4'hF;
    Number1[22][24] = 4'hF;
    Number1[23][24] = 4'hF;
    Number1[0][25] = 4'hF;
    Number1[1][25] = 4'hF;
    Number1[2][25] = 4'hF;
    Number1[3][25] = 4'hF;
    Number1[4][25] = 4'hF;
    Number1[5][25] = 4'hF;
    Number1[6][25] = 4'hF;
    Number1[7][25] = 4'hF;
    Number1[8][25] = 4'hF;
    Number1[9][25] = 4'hF;
    Number1[10][25] = 4'hF;
    Number1[11][25] = 4'hF;
    Number1[12][25] = 4'hC;
    Number1[13][25] = 4'hC;
    Number1[14][25] = 4'hC;
    Number1[15][25] = 4'hC;
    Number1[16][25] = 4'hC;
    Number1[17][25] = 4'hF;
    Number1[18][25] = 4'hF;
    Number1[19][25] = 4'hF;
    Number1[20][25] = 4'hF;
    Number1[21][25] = 4'hF;
    Number1[22][25] = 4'hF;
    Number1[23][25] = 4'hF;
    Number1[0][26] = 4'hF;
    Number1[1][26] = 4'hF;
    Number1[2][26] = 4'hF;
    Number1[3][26] = 4'hF;
    Number1[4][26] = 4'hF;
    Number1[5][26] = 4'hF;
    Number1[6][26] = 4'hF;
    Number1[7][26] = 4'hF;
    Number1[8][26] = 4'hF;
    Number1[9][26] = 4'hF;
    Number1[10][26] = 4'hF;
    Number1[11][26] = 4'hF;
    Number1[12][26] = 4'hC;
    Number1[13][26] = 4'hC;
    Number1[14][26] = 4'hC;
    Number1[15][26] = 4'hC;
    Number1[16][26] = 4'hC;
    Number1[17][26] = 4'hF;
    Number1[18][26] = 4'hF;
    Number1[19][26] = 4'hF;
    Number1[20][26] = 4'hF;
    Number1[21][26] = 4'hF;
    Number1[22][26] = 4'hF;
    Number1[23][26] = 4'hF;
    Number1[0][27] = 4'hF;
    Number1[1][27] = 4'hF;
    Number1[2][27] = 4'hF;
    Number1[3][27] = 4'hF;
    Number1[4][27] = 4'hF;
    Number1[5][27] = 4'hF;
    Number1[6][27] = 4'hF;
    Number1[7][27] = 4'hF;
    Number1[8][27] = 4'hF;
    Number1[9][27] = 4'hF;
    Number1[10][27] = 4'hF;
    Number1[11][27] = 4'hF;
    Number1[12][27] = 4'hC;
    Number1[13][27] = 4'hC;
    Number1[14][27] = 4'hC;
    Number1[15][27] = 4'hC;
    Number1[16][27] = 4'hC;
    Number1[17][27] = 4'hF;
    Number1[18][27] = 4'hF;
    Number1[19][27] = 4'hF;
    Number1[20][27] = 4'hF;
    Number1[21][27] = 4'hF;
    Number1[22][27] = 4'hF;
    Number1[23][27] = 4'hF;
    Number1[0][28] = 4'hF;
    Number1[1][28] = 4'hF;
    Number1[2][28] = 4'hF;
    Number1[3][28] = 4'hF;
    Number1[4][28] = 4'hF;
    Number1[5][28] = 4'hF;
    Number1[6][28] = 4'hF;
    Number1[7][28] = 4'hF;
    Number1[8][28] = 4'hF;
    Number1[9][28] = 4'hF;
    Number1[10][28] = 4'hF;
    Number1[11][28] = 4'hF;
    Number1[12][28] = 4'hF;
    Number1[13][28] = 4'hF;
    Number1[14][28] = 4'hF;
    Number1[15][28] = 4'hF;
    Number1[16][28] = 4'hF;
    Number1[17][28] = 4'hF;
    Number1[18][28] = 4'hF;
    Number1[19][28] = 4'hF;
    Number1[20][28] = 4'hF;
    Number1[21][28] = 4'hF;
    Number1[22][28] = 4'hF;
    Number1[23][28] = 4'hF;
    Number1[0][29] = 4'hF;
    Number1[1][29] = 4'hF;
    Number1[2][29] = 4'hF;
    Number1[3][29] = 4'hF;
    Number1[4][29] = 4'hF;
    Number1[5][29] = 4'hF;
    Number1[6][29] = 4'hF;
    Number1[7][29] = 4'hF;
    Number1[8][29] = 4'hF;
    Number1[9][29] = 4'hF;
    Number1[10][29] = 4'hF;
    Number1[11][29] = 4'hF;
    Number1[12][29] = 4'hF;
    Number1[13][29] = 4'hF;
    Number1[14][29] = 4'hF;
    Number1[15][29] = 4'hF;
    Number1[16][29] = 4'hF;
    Number1[17][29] = 4'hF;
    Number1[18][29] = 4'hF;
    Number1[19][29] = 4'hF;
    Number1[20][29] = 4'hF;
    Number1[21][29] = 4'hF;
    Number1[22][29] = 4'hF;
    Number1[23][29] = 4'hF;
 
//Number 2
    Number2[0][0] = 4'hF;
    Number2[1][0] = 4'hF;
    Number2[2][0] = 4'hF;
    Number2[3][0] = 4'hF;
    Number2[4][0] = 4'hF;
    Number2[5][0] = 4'hF;
    Number2[6][0] = 4'hF;
    Number2[7][0] = 4'hF;
    Number2[8][0] = 4'hF;
    Number2[9][0] = 4'hF;
    Number2[10][0] = 4'hF;
    Number2[11][0] = 4'hF;
    Number2[12][0] = 4'hF;
    Number2[13][0] = 4'hF;
    Number2[14][0] = 4'hF;
    Number2[15][0] = 4'hF;
    Number2[16][0] = 4'hF;
    Number2[17][0] = 4'hF;
    Number2[18][0] = 4'hF;
    Number2[19][0] = 4'hF;
    Number2[20][0] = 4'hF;
    Number2[21][0] = 4'hF;
    Number2[22][0] = 4'hF;
    Number2[23][0] = 4'hF;
    Number2[0][1] = 4'hF;
    Number2[1][1] = 4'hF;
    Number2[2][1] = 4'hF;
    Number2[3][1] = 4'hF;
    Number2[4][1] = 4'hF;
    Number2[5][1] = 4'hF;
    Number2[6][1] = 4'hF;
    Number2[7][1] = 4'hF;
    Number2[8][1] = 4'hF;
    Number2[9][1] = 4'hF;
    Number2[10][1] = 4'hF;
    Number2[11][1] = 4'hF;
    Number2[12][1] = 4'hF;
    Number2[13][1] = 4'hF;
    Number2[14][1] = 4'hF;
    Number2[15][1] = 4'hF;
    Number2[16][1] = 4'hF;
    Number2[17][1] = 4'hF;
    Number2[18][1] = 4'hF;
    Number2[19][1] = 4'hF;
    Number2[20][1] = 4'hF;
    Number2[21][1] = 4'hF;
    Number2[22][1] = 4'hF;
    Number2[23][1] = 4'hF;
    Number2[0][2] = 4'hF;
    Number2[1][2] = 4'hF;
    Number2[2][2] = 4'hF;
    Number2[3][2] = 4'hF;
    Number2[4][2] = 4'hF;
    Number2[5][2] = 4'hF;
    Number2[6][2] = 4'hF;
    Number2[7][2] = 4'hF;
    Number2[8][2] = 4'hF;
    Number2[9][2] = 4'hF;
    Number2[10][2] = 4'hF;
    Number2[11][2] = 4'hF;
    Number2[12][2] = 4'hF;
    Number2[13][2] = 4'hF;
    Number2[14][2] = 4'hF;
    Number2[15][2] = 4'hF;
    Number2[16][2] = 4'hF;
    Number2[17][2] = 4'hF;
    Number2[18][2] = 4'hF;
    Number2[19][2] = 4'hF;
    Number2[20][2] = 4'hF;
    Number2[21][2] = 4'hF;
    Number2[22][2] = 4'hF;
    Number2[23][2] = 4'hF;
    Number2[0][3] = 4'hF;
    Number2[1][3] = 4'hF;
    Number2[2][3] = 4'hC;
    Number2[3][3] = 4'hC;
    Number2[4][3] = 4'hC;
    Number2[5][3] = 4'hC;
    Number2[6][3] = 4'hC;
    Number2[7][3] = 4'hC;
    Number2[8][3] = 4'hC;
    Number2[9][3] = 4'hC;
    Number2[10][3] = 4'hC;
    Number2[11][3] = 4'hC;
    Number2[12][3] = 4'hC;
    Number2[13][3] = 4'hC;
    Number2[14][3] = 4'hC;
    Number2[15][3] = 4'hC;
    Number2[16][3] = 4'hC;
    Number2[17][3] = 4'hF;
    Number2[18][3] = 4'hF;
    Number2[19][3] = 4'hF;
    Number2[20][3] = 4'hF;
    Number2[21][3] = 4'hF;
    Number2[22][3] = 4'hF;
    Number2[23][3] = 4'hF;
    Number2[0][4] = 4'hF;
    Number2[1][4] = 4'hF;
    Number2[2][4] = 4'hC;
    Number2[3][4] = 4'hC;
    Number2[4][4] = 4'hC;
    Number2[5][4] = 4'hC;
    Number2[6][4] = 4'hC;
    Number2[7][4] = 4'hC;
    Number2[8][4] = 4'hC;
    Number2[9][4] = 4'hC;
    Number2[10][4] = 4'hC;
    Number2[11][4] = 4'hC;
    Number2[12][4] = 4'hC;
    Number2[13][4] = 4'hC;
    Number2[14][4] = 4'hC;
    Number2[15][4] = 4'hC;
    Number2[16][4] = 4'hC;
    Number2[17][4] = 4'hF;
    Number2[18][4] = 4'hF;
    Number2[19][4] = 4'hF;
    Number2[20][4] = 4'hF;
    Number2[21][4] = 4'hF;
    Number2[22][4] = 4'hF;
    Number2[23][4] = 4'hF;
    Number2[0][5] = 4'hF;
    Number2[1][5] = 4'hF;
    Number2[2][5] = 4'hC;
    Number2[3][5] = 4'hC;
    Number2[4][5] = 4'hC;
    Number2[5][5] = 4'hC;
    Number2[6][5] = 4'hC;
    Number2[7][5] = 4'hC;
    Number2[8][5] = 4'hC;
    Number2[9][5] = 4'hC;
    Number2[10][5] = 4'hC;
    Number2[11][5] = 4'hC;
    Number2[12][5] = 4'hC;
    Number2[13][5] = 4'hC;
    Number2[14][5] = 4'hC;
    Number2[15][5] = 4'hC;
    Number2[16][5] = 4'hC;
    Number2[17][5] = 4'hF;
    Number2[18][5] = 4'hF;
    Number2[19][5] = 4'hF;
    Number2[20][5] = 4'hF;
    Number2[21][5] = 4'hF;
    Number2[22][5] = 4'hF;
    Number2[23][5] = 4'hF;
    Number2[0][6] = 4'hF;
    Number2[1][6] = 4'hF;
    Number2[2][6] = 4'hC;
    Number2[3][6] = 4'hC;
    Number2[4][6] = 4'hC;
    Number2[5][6] = 4'hC;
    Number2[6][6] = 4'hC;
    Number2[7][6] = 4'hC;
    Number2[8][6] = 4'hC;
    Number2[9][6] = 4'hC;
    Number2[10][6] = 4'hC;
    Number2[11][6] = 4'hC;
    Number2[12][6] = 4'hC;
    Number2[13][6] = 4'hC;
    Number2[14][6] = 4'hC;
    Number2[15][6] = 4'hC;
    Number2[16][6] = 4'hC;
    Number2[17][6] = 4'hF;
    Number2[18][6] = 4'hF;
    Number2[19][6] = 4'hF;
    Number2[20][6] = 4'hF;
    Number2[21][6] = 4'hF;
    Number2[22][6] = 4'hF;
    Number2[23][6] = 4'hF;
    Number2[0][7] = 4'hF;
    Number2[1][7] = 4'hF;
    Number2[2][7] = 4'hC;
    Number2[3][7] = 4'hC;
    Number2[4][7] = 4'hC;
    Number2[5][7] = 4'hC;
    Number2[6][7] = 4'hC;
    Number2[7][7] = 4'hC;
    Number2[8][7] = 4'hC;
    Number2[9][7] = 4'hC;
    Number2[10][7] = 4'hC;
    Number2[11][7] = 4'hC;
    Number2[12][7] = 4'hC;
    Number2[13][7] = 4'hC;
    Number2[14][7] = 4'hC;
    Number2[15][7] = 4'hC;
    Number2[16][7] = 4'hC;
    Number2[17][7] = 4'hF;
    Number2[18][7] = 4'hF;
    Number2[19][7] = 4'hF;
    Number2[20][7] = 4'hF;
    Number2[21][7] = 4'hF;
    Number2[22][7] = 4'hF;
    Number2[23][7] = 4'hF;
    Number2[0][8] = 4'hF;
    Number2[1][8] = 4'hF;
    Number2[2][8] = 4'hF;
    Number2[3][8] = 4'hF;
    Number2[4][8] = 4'hF;
    Number2[5][8] = 4'hF;
    Number2[6][8] = 4'hF;
    Number2[7][8] = 4'hF;
    Number2[8][8] = 4'hF;
    Number2[9][8] = 4'hF;
    Number2[10][8] = 4'hF;
    Number2[11][8] = 4'hF;
    Number2[12][8] = 4'hF;
    Number2[13][8] = 4'hF;
    Number2[14][8] = 4'hF;
    Number2[15][8] = 4'hF;
    Number2[16][8] = 4'hF;
    Number2[17][8] = 4'hC;
    Number2[18][8] = 4'hC;
    Number2[19][8] = 4'hC;
    Number2[20][8] = 4'hC;
    Number2[21][8] = 4'hC;
    Number2[22][8] = 4'hF;
    Number2[23][8] = 4'hF;
    Number2[0][9] = 4'hF;
    Number2[1][9] = 4'hF;
    Number2[2][9] = 4'hF;
    Number2[3][9] = 4'hF;
    Number2[4][9] = 4'hF;
    Number2[5][9] = 4'hF;
    Number2[6][9] = 4'hF;
    Number2[7][9] = 4'hF;
    Number2[8][9] = 4'hF;
    Number2[9][9] = 4'hF;
    Number2[10][9] = 4'hF;
    Number2[11][9] = 4'hF;
    Number2[12][9] = 4'hF;
    Number2[13][9] = 4'hF;
    Number2[14][9] = 4'hF;
    Number2[15][9] = 4'hF;
    Number2[16][9] = 4'hF;
    Number2[17][9] = 4'hC;
    Number2[18][9] = 4'hC;
    Number2[19][9] = 4'hC;
    Number2[20][9] = 4'hC;
    Number2[21][9] = 4'hC;
    Number2[22][9] = 4'hF;
    Number2[23][9] = 4'hF;
    Number2[0][10] = 4'hF;
    Number2[1][10] = 4'hF;
    Number2[2][10] = 4'hF;
    Number2[3][10] = 4'hF;
    Number2[4][10] = 4'hF;
    Number2[5][10] = 4'hF;
    Number2[6][10] = 4'hF;
    Number2[7][10] = 4'hF;
    Number2[8][10] = 4'hF;
    Number2[9][10] = 4'hF;
    Number2[10][10] = 4'hF;
    Number2[11][10] = 4'hF;
    Number2[12][10] = 4'hF;
    Number2[13][10] = 4'hF;
    Number2[14][10] = 4'hF;
    Number2[15][10] = 4'hF;
    Number2[16][10] = 4'hF;
    Number2[17][10] = 4'hC;
    Number2[18][10] = 4'hC;
    Number2[19][10] = 4'hC;
    Number2[20][10] = 4'hC;
    Number2[21][10] = 4'hC;
    Number2[22][10] = 4'hF;
    Number2[23][10] = 4'hF;
    Number2[0][11] = 4'hF;
    Number2[1][11] = 4'hF;
    Number2[2][11] = 4'hF;
    Number2[3][11] = 4'hF;
    Number2[4][11] = 4'hF;
    Number2[5][11] = 4'hF;
    Number2[6][11] = 4'hF;
    Number2[7][11] = 4'hF;
    Number2[8][11] = 4'hF;
    Number2[9][11] = 4'hF;
    Number2[10][11] = 4'hF;
    Number2[11][11] = 4'hF;
    Number2[12][11] = 4'hF;
    Number2[13][11] = 4'hF;
    Number2[14][11] = 4'hF;
    Number2[15][11] = 4'hF;
    Number2[16][11] = 4'hF;
    Number2[17][11] = 4'hC;
    Number2[18][11] = 4'hC;
    Number2[19][11] = 4'hC;
    Number2[20][11] = 4'hC;
    Number2[21][11] = 4'hC;
    Number2[22][11] = 4'hF;
    Number2[23][11] = 4'hF;
    Number2[0][12] = 4'hF;
    Number2[1][12] = 4'hF;
    Number2[2][12] = 4'hF;
    Number2[3][12] = 4'hF;
    Number2[4][12] = 4'hF;
    Number2[5][12] = 4'hF;
    Number2[6][12] = 4'hF;
    Number2[7][12] = 4'hF;
    Number2[8][12] = 4'hF;
    Number2[9][12] = 4'hF;
    Number2[10][12] = 4'hF;
    Number2[11][12] = 4'hF;
    Number2[12][12] = 4'hF;
    Number2[13][12] = 4'hF;
    Number2[14][12] = 4'hF;
    Number2[15][12] = 4'hF;
    Number2[16][12] = 4'hF;
    Number2[17][12] = 4'hC;
    Number2[18][12] = 4'hC;
    Number2[19][12] = 4'hC;
    Number2[20][12] = 4'hC;
    Number2[21][12] = 4'hC;
    Number2[22][12] = 4'hF;
    Number2[23][12] = 4'hF;
    Number2[0][13] = 4'hF;
    Number2[1][13] = 4'hF;
    Number2[2][13] = 4'hF;
    Number2[3][13] = 4'hF;
    Number2[4][13] = 4'hF;
    Number2[5][13] = 4'hF;
    Number2[6][13] = 4'hF;
    Number2[7][13] = 4'hC;
    Number2[8][13] = 4'hC;
    Number2[9][13] = 4'hC;
    Number2[10][13] = 4'hC;
    Number2[11][13] = 4'hC;
    Number2[12][13] = 4'hC;
    Number2[13][13] = 4'hC;
    Number2[14][13] = 4'hC;
    Number2[15][13] = 4'hC;
    Number2[16][13] = 4'hC;
    Number2[17][13] = 4'hF;
    Number2[18][13] = 4'hF;
    Number2[19][13] = 4'hF;
    Number2[20][13] = 4'hF;
    Number2[21][13] = 4'hF;
    Number2[22][13] = 4'hF;
    Number2[23][13] = 4'hF;
    Number2[0][14] = 4'hF;
    Number2[1][14] = 4'hF;
    Number2[2][14] = 4'hF;
    Number2[3][14] = 4'hF;
    Number2[4][14] = 4'hF;
    Number2[5][14] = 4'hF;
    Number2[6][14] = 4'hF;
    Number2[7][14] = 4'hC;
    Number2[8][14] = 4'hC;
    Number2[9][14] = 4'hC;
    Number2[10][14] = 4'hC;
    Number2[11][14] = 4'hC;
    Number2[12][14] = 4'hC;
    Number2[13][14] = 4'hC;
    Number2[14][14] = 4'hC;
    Number2[15][14] = 4'hC;
    Number2[16][14] = 4'hC;
    Number2[17][14] = 4'hF;
    Number2[18][14] = 4'hF;
    Number2[19][14] = 4'hF;
    Number2[20][14] = 4'hF;
    Number2[21][14] = 4'hF;
    Number2[22][14] = 4'hF;
    Number2[23][14] = 4'hF;
    Number2[0][15] = 4'hF;
    Number2[1][15] = 4'hF;
    Number2[2][15] = 4'hF;
    Number2[3][15] = 4'hF;
    Number2[4][15] = 4'hF;
    Number2[5][15] = 4'hF;
    Number2[6][15] = 4'hF;
    Number2[7][15] = 4'hC;
    Number2[8][15] = 4'hC;
    Number2[9][15] = 4'hC;
    Number2[10][15] = 4'hC;
    Number2[11][15] = 4'hC;
    Number2[12][15] = 4'hC;
    Number2[13][15] = 4'hC;
    Number2[14][15] = 4'hC;
    Number2[15][15] = 4'hC;
    Number2[16][15] = 4'hC;
    Number2[17][15] = 4'hF;
    Number2[18][15] = 4'hF;
    Number2[19][15] = 4'hF;
    Number2[20][15] = 4'hF;
    Number2[21][15] = 4'hF;
    Number2[22][15] = 4'hF;
    Number2[23][15] = 4'hF;
    Number2[0][16] = 4'hF;
    Number2[1][16] = 4'hF;
    Number2[2][16] = 4'hF;
    Number2[3][16] = 4'hF;
    Number2[4][16] = 4'hF;
    Number2[5][16] = 4'hF;
    Number2[6][16] = 4'hF;
    Number2[7][16] = 4'hC;
    Number2[8][16] = 4'hC;
    Number2[9][16] = 4'hC;
    Number2[10][16] = 4'hC;
    Number2[11][16] = 4'hC;
    Number2[12][16] = 4'hC;
    Number2[13][16] = 4'hC;
    Number2[14][16] = 4'hC;
    Number2[15][16] = 4'hC;
    Number2[16][16] = 4'hC;
    Number2[17][16] = 4'hF;
    Number2[18][16] = 4'hF;
    Number2[19][16] = 4'hF;
    Number2[20][16] = 4'hF;
    Number2[21][16] = 4'hF;
    Number2[22][16] = 4'hF;
    Number2[23][16] = 4'hF;
    Number2[0][17] = 4'hF;
    Number2[1][17] = 4'hF;
    Number2[2][17] = 4'hF;
    Number2[3][17] = 4'hF;
    Number2[4][17] = 4'hF;
    Number2[5][17] = 4'hF;
    Number2[6][17] = 4'hF;
    Number2[7][17] = 4'hC;
    Number2[8][17] = 4'hC;
    Number2[9][17] = 4'hC;
    Number2[10][17] = 4'hC;
    Number2[11][17] = 4'hC;
    Number2[12][17] = 4'hC;
    Number2[13][17] = 4'hC;
    Number2[14][17] = 4'hC;
    Number2[15][17] = 4'hC;
    Number2[16][17] = 4'hC;
    Number2[17][17] = 4'hF;
    Number2[18][17] = 4'hF;
    Number2[19][17] = 4'hF;
    Number2[20][17] = 4'hF;
    Number2[21][17] = 4'hF;
    Number2[22][17] = 4'hF;
    Number2[23][17] = 4'hF;
    Number2[0][18] = 4'hF;
    Number2[1][18] = 4'hF;
    Number2[2][18] = 4'hC;
    Number2[3][18] = 4'hC;
    Number2[4][18] = 4'hC;
    Number2[5][18] = 4'hC;
    Number2[6][18] = 4'hC;
    Number2[7][18] = 4'hF;
    Number2[8][18] = 4'hF;
    Number2[9][18] = 4'hF;
    Number2[10][18] = 4'hF;
    Number2[11][18] = 4'hF;
    Number2[12][18] = 4'hF;
    Number2[13][18] = 4'hF;
    Number2[14][18] = 4'hF;
    Number2[15][18] = 4'hF;
    Number2[16][18] = 4'hF;
    Number2[17][18] = 4'hF;
    Number2[18][18] = 4'hF;
    Number2[19][18] = 4'hF;
    Number2[20][18] = 4'hF;
    Number2[21][18] = 4'hF;
    Number2[22][18] = 4'hF;
    Number2[23][18] = 4'hF;
    Number2[0][19] = 4'hF;
    Number2[1][19] = 4'hF;
    Number2[2][19] = 4'hC;
    Number2[3][19] = 4'hC;
    Number2[4][19] = 4'hC;
    Number2[5][19] = 4'hC;
    Number2[6][19] = 4'hC;
    Number2[7][19] = 4'hF;
    Number2[8][19] = 4'hF;
    Number2[9][19] = 4'hF;
    Number2[10][19] = 4'hF;
    Number2[11][19] = 4'hF;
    Number2[12][19] = 4'hF;
    Number2[13][19] = 4'hF;
    Number2[14][19] = 4'hF;
    Number2[15][19] = 4'hF;
    Number2[16][19] = 4'hF;
    Number2[17][19] = 4'hF;
    Number2[18][19] = 4'hF;
    Number2[19][19] = 4'hF;
    Number2[20][19] = 4'hF;
    Number2[21][19] = 4'hF;
    Number2[22][19] = 4'hF;
    Number2[23][19] = 4'hF;
    Number2[0][20] = 4'hF;
    Number2[1][20] = 4'hF;
    Number2[2][20] = 4'hC;
    Number2[3][20] = 4'hC;
    Number2[4][20] = 4'hC;
    Number2[5][20] = 4'hC;
    Number2[6][20] = 4'hC;
    Number2[7][20] = 4'hF;
    Number2[8][20] = 4'hF;
    Number2[9][20] = 4'hF;
    Number2[10][20] = 4'hF;
    Number2[11][20] = 4'hF;
    Number2[12][20] = 4'hF;
    Number2[13][20] = 4'hF;
    Number2[14][20] = 4'hF;
    Number2[15][20] = 4'hF;
    Number2[16][20] = 4'hF;
    Number2[17][20] = 4'hF;
    Number2[18][20] = 4'hF;
    Number2[19][20] = 4'hF;
    Number2[20][20] = 4'hF;
    Number2[21][20] = 4'hF;
    Number2[22][20] = 4'hF;
    Number2[23][20] = 4'hF;
    Number2[0][21] = 4'hF;
    Number2[1][21] = 4'hF;
    Number2[2][21] = 4'hC;
    Number2[3][21] = 4'hC;
    Number2[4][21] = 4'hC;
    Number2[5][21] = 4'hC;
    Number2[6][21] = 4'hC;
    Number2[7][21] = 4'hF;
    Number2[8][21] = 4'hF;
    Number2[9][21] = 4'hF;
    Number2[10][21] = 4'hF;
    Number2[11][21] = 4'hF;
    Number2[12][21] = 4'hF;
    Number2[13][21] = 4'hF;
    Number2[14][21] = 4'hF;
    Number2[15][21] = 4'hF;
    Number2[16][21] = 4'hF;
    Number2[17][21] = 4'hF;
    Number2[18][21] = 4'hF;
    Number2[19][21] = 4'hF;
    Number2[20][21] = 4'hF;
    Number2[21][21] = 4'hF;
    Number2[22][21] = 4'hF;
    Number2[23][21] = 4'hF;
    Number2[0][22] = 4'hF;
    Number2[1][22] = 4'hF;
    Number2[2][22] = 4'hC;
    Number2[3][22] = 4'hC;
    Number2[4][22] = 4'hC;
    Number2[5][22] = 4'hC;
    Number2[6][22] = 4'hC;
    Number2[7][22] = 4'hF;
    Number2[8][22] = 4'hF;
    Number2[9][22] = 4'hF;
    Number2[10][22] = 4'hF;
    Number2[11][22] = 4'hF;
    Number2[12][22] = 4'hF;
    Number2[13][22] = 4'hF;
    Number2[14][22] = 4'hF;
    Number2[15][22] = 4'hF;
    Number2[16][22] = 4'hF;
    Number2[17][22] = 4'hF;
    Number2[18][22] = 4'hF;
    Number2[19][22] = 4'hF;
    Number2[20][22] = 4'hF;
    Number2[21][22] = 4'hF;
    Number2[22][22] = 4'hF;
    Number2[23][22] = 4'hF;
    Number2[0][23] = 4'hF;
    Number2[1][23] = 4'hF;
    Number2[2][23] = 4'hC;
    Number2[3][23] = 4'hC;
    Number2[4][23] = 4'hC;
    Number2[5][23] = 4'hC;
    Number2[6][23] = 4'hC;
    Number2[7][23] = 4'hC;
    Number2[8][23] = 4'hC;
    Number2[9][23] = 4'hC;
    Number2[10][23] = 4'hC;
    Number2[11][23] = 4'hC;
    Number2[12][23] = 4'hC;
    Number2[13][23] = 4'hC;
    Number2[14][23] = 4'hC;
    Number2[15][23] = 4'hC;
    Number2[16][23] = 4'hC;
    Number2[17][23] = 4'hC;
    Number2[18][23] = 4'hC;
    Number2[19][23] = 4'hC;
    Number2[20][23] = 4'hC;
    Number2[21][23] = 4'hC;
    Number2[22][23] = 4'hF;
    Number2[23][23] = 4'hF;
    Number2[0][24] = 4'hF;
    Number2[1][24] = 4'hF;
    Number2[2][24] = 4'hC;
    Number2[3][24] = 4'hC;
    Number2[4][24] = 4'hC;
    Number2[5][24] = 4'hC;
    Number2[6][24] = 4'hC;
    Number2[7][24] = 4'hC;
    Number2[8][24] = 4'hC;
    Number2[9][24] = 4'hC;
    Number2[10][24] = 4'hC;
    Number2[11][24] = 4'hC;
    Number2[12][24] = 4'hC;
    Number2[13][24] = 4'hC;
    Number2[14][24] = 4'hC;
    Number2[15][24] = 4'hC;
    Number2[16][24] = 4'hC;
    Number2[17][24] = 4'hC;
    Number2[18][24] = 4'hC;
    Number2[19][24] = 4'hC;
    Number2[20][24] = 4'hC;
    Number2[21][24] = 4'hC;
    Number2[22][24] = 4'hF;
    Number2[23][24] = 4'hF;
    Number2[0][25] = 4'hF;
    Number2[1][25] = 4'hF;
    Number2[2][25] = 4'hC;
    Number2[3][25] = 4'hC;
    Number2[4][25] = 4'hC;
    Number2[5][25] = 4'hC;
    Number2[6][25] = 4'hC;
    Number2[7][25] = 4'hC;
    Number2[8][25] = 4'hC;
    Number2[9][25] = 4'hC;
    Number2[10][25] = 4'hC;
    Number2[11][25] = 4'hC;
    Number2[12][25] = 4'hC;
    Number2[13][25] = 4'hC;
    Number2[14][25] = 4'hC;
    Number2[15][25] = 4'hC;
    Number2[16][25] = 4'hC;
    Number2[17][25] = 4'hC;
    Number2[18][25] = 4'hC;
    Number2[19][25] = 4'hC;
    Number2[20][25] = 4'hC;
    Number2[21][25] = 4'hC;
    Number2[22][25] = 4'hF;
    Number2[23][25] = 4'hF;
    Number2[0][26] = 4'hF;
    Number2[1][26] = 4'hF;
    Number2[2][26] = 4'hC;
    Number2[3][26] = 4'hC;
    Number2[4][26] = 4'hC;
    Number2[5][26] = 4'hC;
    Number2[6][26] = 4'hC;
    Number2[7][26] = 4'hC;
    Number2[8][26] = 4'hC;
    Number2[9][26] = 4'hC;
    Number2[10][26] = 4'hC;
    Number2[11][26] = 4'hC;
    Number2[12][26] = 4'hC;
    Number2[13][26] = 4'hC;
    Number2[14][26] = 4'hC;
    Number2[15][26] = 4'hC;
    Number2[16][26] = 4'hC;
    Number2[17][26] = 4'hC;
    Number2[18][26] = 4'hC;
    Number2[19][26] = 4'hC;
    Number2[20][26] = 4'hC;
    Number2[21][26] = 4'hC;
    Number2[22][26] = 4'hF;
    Number2[23][26] = 4'hF;
    Number2[0][27] = 4'hF;
    Number2[1][27] = 4'hF;
    Number2[2][27] = 4'hC;
    Number2[3][27] = 4'hC;
    Number2[4][27] = 4'hC;
    Number2[5][27] = 4'hC;
    Number2[6][27] = 4'hC;
    Number2[7][27] = 4'hC;
    Number2[8][27] = 4'hC;
    Number2[9][27] = 4'hC;
    Number2[10][27] = 4'hC;
    Number2[11][27] = 4'hC;
    Number2[12][27] = 4'hC;
    Number2[13][27] = 4'hC;
    Number2[14][27] = 4'hC;
    Number2[15][27] = 4'hC;
    Number2[16][27] = 4'hC;
    Number2[17][27] = 4'hC;
    Number2[18][27] = 4'hC;
    Number2[19][27] = 4'hC;
    Number2[20][27] = 4'hC;
    Number2[21][27] = 4'hC;
    Number2[22][27] = 4'hF;
    Number2[23][27] = 4'hF;
    Number2[0][28] = 4'hF;
    Number2[1][28] = 4'hF;
    Number2[2][28] = 4'hF;
    Number2[3][28] = 4'hF;
    Number2[4][28] = 4'hF;
    Number2[5][28] = 4'hF;
    Number2[6][28] = 4'hF;
    Number2[7][28] = 4'hF;
    Number2[8][28] = 4'hF;
    Number2[9][28] = 4'hF;
    Number2[10][28] = 4'hF;
    Number2[11][28] = 4'hF;
    Number2[12][28] = 4'hF;
    Number2[13][28] = 4'hF;
    Number2[14][28] = 4'hF;
    Number2[15][28] = 4'hF;
    Number2[16][28] = 4'hF;
    Number2[17][28] = 4'hF;
    Number2[18][28] = 4'hF;
    Number2[19][28] = 4'hF;
    Number2[20][28] = 4'hF;
    Number2[21][28] = 4'hF;
    Number2[22][28] = 4'hF;
    Number2[23][28] = 4'hF;
    Number2[0][29] = 4'hF;
    Number2[1][29] = 4'hF;
    Number2[2][29] = 4'hF;
    Number2[3][29] = 4'hF;
    Number2[4][29] = 4'hF;
    Number2[5][29] = 4'hF;
    Number2[6][29] = 4'hF;
    Number2[7][29] = 4'hF;
    Number2[8][29] = 4'hF;
    Number2[9][29] = 4'hF;
    Number2[10][29] = 4'hF;
    Number2[11][29] = 4'hF;
    Number2[12][29] = 4'hF;
    Number2[13][29] = 4'hF;
    Number2[14][29] = 4'hF;
    Number2[15][29] = 4'hF;
    Number2[16][29] = 4'hF;
    Number2[17][29] = 4'hF;
    Number2[18][29] = 4'hF;
    Number2[19][29] = 4'hF;
    Number2[20][29] = 4'hF;
    Number2[21][29] = 4'hF;
    Number2[22][29] = 4'hF;
    Number2[23][29] = 4'hF;
 
//Number 3
    Number3[0][0] = 4'hF;
    Number3[1][0] = 4'hF;
    Number3[2][0] = 4'hF;
    Number3[3][0] = 4'hF;
    Number3[4][0] = 4'hF;
    Number3[5][0] = 4'hF;
    Number3[6][0] = 4'hF;
    Number3[7][0] = 4'hF;
    Number3[8][0] = 4'hF;
    Number3[9][0] = 4'hF;
    Number3[10][0] = 4'hF;
    Number3[11][0] = 4'hF;
    Number3[12][0] = 4'hF;
    Number3[13][0] = 4'hF;
    Number3[14][0] = 4'hF;
    Number3[15][0] = 4'hF;
    Number3[16][0] = 4'hF;
    Number3[17][0] = 4'hF;
    Number3[18][0] = 4'hF;
    Number3[19][0] = 4'hF;
    Number3[20][0] = 4'hF;
    Number3[21][0] = 4'hF;
    Number3[22][0] = 4'hF;
    Number3[23][0] = 4'hF;
    Number3[0][1] = 4'hF;
    Number3[1][1] = 4'hF;
    Number3[2][1] = 4'hF;
    Number3[3][1] = 4'hF;
    Number3[4][1] = 4'hF;
    Number3[5][1] = 4'hF;
    Number3[6][1] = 4'hF;
    Number3[7][1] = 4'hF;
    Number3[8][1] = 4'hF;
    Number3[9][1] = 4'hF;
    Number3[10][1] = 4'hF;
    Number3[11][1] = 4'hF;
    Number3[12][1] = 4'hF;
    Number3[13][1] = 4'hF;
    Number3[14][1] = 4'hF;
    Number3[15][1] = 4'hF;
    Number3[16][1] = 4'hF;
    Number3[17][1] = 4'hF;
    Number3[18][1] = 4'hF;
    Number3[19][1] = 4'hF;
    Number3[20][1] = 4'hF;
    Number3[21][1] = 4'hF;
    Number3[22][1] = 4'hF;
    Number3[23][1] = 4'hF;
    Number3[0][2] = 4'hF;
    Number3[1][2] = 4'hF;
    Number3[2][2] = 4'hF;
    Number3[3][2] = 4'hF;
    Number3[4][2] = 4'hF;
    Number3[5][2] = 4'hF;
    Number3[6][2] = 4'hF;
    Number3[7][2] = 4'hF;
    Number3[8][2] = 4'hF;
    Number3[9][2] = 4'hF;
    Number3[10][2] = 4'hF;
    Number3[11][2] = 4'hF;
    Number3[12][2] = 4'hF;
    Number3[13][2] = 4'hF;
    Number3[14][2] = 4'hF;
    Number3[15][2] = 4'hF;
    Number3[16][2] = 4'hF;
    Number3[17][2] = 4'hF;
    Number3[18][2] = 4'hF;
    Number3[19][2] = 4'hF;
    Number3[20][2] = 4'hF;
    Number3[21][2] = 4'hF;
    Number3[22][2] = 4'hF;
    Number3[23][2] = 4'hF;
    Number3[0][3] = 4'hF;
    Number3[1][3] = 4'hF;
    Number3[2][3] = 4'hC;
    Number3[3][3] = 4'hC;
    Number3[4][3] = 4'hC;
    Number3[5][3] = 4'hC;
    Number3[6][3] = 4'hC;
    Number3[7][3] = 4'hC;
    Number3[8][3] = 4'hC;
    Number3[9][3] = 4'hC;
    Number3[10][3] = 4'hC;
    Number3[11][3] = 4'hC;
    Number3[12][3] = 4'hC;
    Number3[13][3] = 4'hC;
    Number3[14][3] = 4'hC;
    Number3[15][3] = 4'hC;
    Number3[16][3] = 4'hC;
    Number3[17][3] = 4'hF;
    Number3[18][3] = 4'hF;
    Number3[19][3] = 4'hF;
    Number3[20][3] = 4'hF;
    Number3[21][3] = 4'hF;
    Number3[22][3] = 4'hF;
    Number3[23][3] = 4'hF;
    Number3[0][4] = 4'hF;
    Number3[1][4] = 4'hF;
    Number3[2][4] = 4'hC;
    Number3[3][4] = 4'hC;
    Number3[4][4] = 4'hC;
    Number3[5][4] = 4'hC;
    Number3[6][4] = 4'hC;
    Number3[7][4] = 4'hC;
    Number3[8][4] = 4'hC;
    Number3[9][4] = 4'hC;
    Number3[10][4] = 4'hC;
    Number3[11][4] = 4'hC;
    Number3[12][4] = 4'hC;
    Number3[13][4] = 4'hC;
    Number3[14][4] = 4'hC;
    Number3[15][4] = 4'hC;
    Number3[16][4] = 4'hC;
    Number3[17][4] = 4'hF;
    Number3[18][4] = 4'hF;
    Number3[19][4] = 4'hF;
    Number3[20][4] = 4'hF;
    Number3[21][4] = 4'hF;
    Number3[22][4] = 4'hF;
    Number3[23][4] = 4'hF;
    Number3[0][5] = 4'hF;
    Number3[1][5] = 4'hF;
    Number3[2][5] = 4'hC;
    Number3[3][5] = 4'hC;
    Number3[4][5] = 4'hC;
    Number3[5][5] = 4'hC;
    Number3[6][5] = 4'hC;
    Number3[7][5] = 4'hC;
    Number3[8][5] = 4'hC;
    Number3[9][5] = 4'hC;
    Number3[10][5] = 4'hC;
    Number3[11][5] = 4'hC;
    Number3[12][5] = 4'hC;
    Number3[13][5] = 4'hC;
    Number3[14][5] = 4'hC;
    Number3[15][5] = 4'hC;
    Number3[16][5] = 4'hC;
    Number3[17][5] = 4'hF;
    Number3[18][5] = 4'hF;
    Number3[19][5] = 4'hF;
    Number3[20][5] = 4'hF;
    Number3[21][5] = 4'hF;
    Number3[22][5] = 4'hF;
    Number3[23][5] = 4'hF;
    Number3[0][6] = 4'hF;
    Number3[1][6] = 4'hF;
    Number3[2][6] = 4'hC;
    Number3[3][6] = 4'hC;
    Number3[4][6] = 4'hC;
    Number3[5][6] = 4'hC;
    Number3[6][6] = 4'hC;
    Number3[7][6] = 4'hC;
    Number3[8][6] = 4'hC;
    Number3[9][6] = 4'hC;
    Number3[10][6] = 4'hC;
    Number3[11][6] = 4'hC;
    Number3[12][6] = 4'hC;
    Number3[13][6] = 4'hC;
    Number3[14][6] = 4'hC;
    Number3[15][6] = 4'hC;
    Number3[16][6] = 4'hC;
    Number3[17][6] = 4'hF;
    Number3[18][6] = 4'hF;
    Number3[19][6] = 4'hF;
    Number3[20][6] = 4'hF;
    Number3[21][6] = 4'hF;
    Number3[22][6] = 4'hF;
    Number3[23][6] = 4'hF;
    Number3[0][7] = 4'hF;
    Number3[1][7] = 4'hF;
    Number3[2][7] = 4'hC;
    Number3[3][7] = 4'hC;
    Number3[4][7] = 4'hC;
    Number3[5][7] = 4'hC;
    Number3[6][7] = 4'hC;
    Number3[7][7] = 4'hC;
    Number3[8][7] = 4'hC;
    Number3[9][7] = 4'hC;
    Number3[10][7] = 4'hC;
    Number3[11][7] = 4'hC;
    Number3[12][7] = 4'hC;
    Number3[13][7] = 4'hC;
    Number3[14][7] = 4'hC;
    Number3[15][7] = 4'hC;
    Number3[16][7] = 4'hC;
    Number3[17][7] = 4'hF;
    Number3[18][7] = 4'hF;
    Number3[19][7] = 4'hF;
    Number3[20][7] = 4'hF;
    Number3[21][7] = 4'hF;
    Number3[22][7] = 4'hF;
    Number3[23][7] = 4'hF;
    Number3[0][8] = 4'hF;
    Number3[1][8] = 4'hF;
    Number3[2][8] = 4'hF;
    Number3[3][8] = 4'hF;
    Number3[4][8] = 4'hF;
    Number3[5][8] = 4'hF;
    Number3[6][8] = 4'hF;
    Number3[7][8] = 4'hF;
    Number3[8][8] = 4'hF;
    Number3[9][8] = 4'hF;
    Number3[10][8] = 4'hF;
    Number3[11][8] = 4'hF;
    Number3[12][8] = 4'hF;
    Number3[13][8] = 4'hF;
    Number3[14][8] = 4'hF;
    Number3[15][8] = 4'hF;
    Number3[16][8] = 4'hF;
    Number3[17][8] = 4'hC;
    Number3[18][8] = 4'hC;
    Number3[19][8] = 4'hC;
    Number3[20][8] = 4'hC;
    Number3[21][8] = 4'hC;
    Number3[22][8] = 4'hF;
    Number3[23][8] = 4'hF;
    Number3[0][9] = 4'hF;
    Number3[1][9] = 4'hF;
    Number3[2][9] = 4'hF;
    Number3[3][9] = 4'hF;
    Number3[4][9] = 4'hF;
    Number3[5][9] = 4'hF;
    Number3[6][9] = 4'hF;
    Number3[7][9] = 4'hF;
    Number3[8][9] = 4'hF;
    Number3[9][9] = 4'hF;
    Number3[10][9] = 4'hF;
    Number3[11][9] = 4'hF;
    Number3[12][9] = 4'hF;
    Number3[13][9] = 4'hF;
    Number3[14][9] = 4'hF;
    Number3[15][9] = 4'hF;
    Number3[16][9] = 4'hF;
    Number3[17][9] = 4'hC;
    Number3[18][9] = 4'hC;
    Number3[19][9] = 4'hC;
    Number3[20][9] = 4'hC;
    Number3[21][9] = 4'hC;
    Number3[22][9] = 4'hF;
    Number3[23][9] = 4'hF;
    Number3[0][10] = 4'hF;
    Number3[1][10] = 4'hF;
    Number3[2][10] = 4'hF;
    Number3[3][10] = 4'hF;
    Number3[4][10] = 4'hF;
    Number3[5][10] = 4'hF;
    Number3[6][10] = 4'hF;
    Number3[7][10] = 4'hF;
    Number3[8][10] = 4'hF;
    Number3[9][10] = 4'hF;
    Number3[10][10] = 4'hF;
    Number3[11][10] = 4'hF;
    Number3[12][10] = 4'hF;
    Number3[13][10] = 4'hF;
    Number3[14][10] = 4'hF;
    Number3[15][10] = 4'hF;
    Number3[16][10] = 4'hF;
    Number3[17][10] = 4'hC;
    Number3[18][10] = 4'hC;
    Number3[19][10] = 4'hC;
    Number3[20][10] = 4'hC;
    Number3[21][10] = 4'hC;
    Number3[22][10] = 4'hF;
    Number3[23][10] = 4'hF;
    Number3[0][11] = 4'hF;
    Number3[1][11] = 4'hF;
    Number3[2][11] = 4'hF;
    Number3[3][11] = 4'hF;
    Number3[4][11] = 4'hF;
    Number3[5][11] = 4'hF;
    Number3[6][11] = 4'hF;
    Number3[7][11] = 4'hF;
    Number3[8][11] = 4'hF;
    Number3[9][11] = 4'hF;
    Number3[10][11] = 4'hF;
    Number3[11][11] = 4'hF;
    Number3[12][11] = 4'hF;
    Number3[13][11] = 4'hF;
    Number3[14][11] = 4'hF;
    Number3[15][11] = 4'hF;
    Number3[16][11] = 4'hF;
    Number3[17][11] = 4'hC;
    Number3[18][11] = 4'hC;
    Number3[19][11] = 4'hC;
    Number3[20][11] = 4'hC;
    Number3[21][11] = 4'hC;
    Number3[22][11] = 4'hF;
    Number3[23][11] = 4'hF;
    Number3[0][12] = 4'hF;
    Number3[1][12] = 4'hF;
    Number3[2][12] = 4'hF;
    Number3[3][12] = 4'hF;
    Number3[4][12] = 4'hF;
    Number3[5][12] = 4'hF;
    Number3[6][12] = 4'hF;
    Number3[7][12] = 4'hF;
    Number3[8][12] = 4'hF;
    Number3[9][12] = 4'hF;
    Number3[10][12] = 4'hF;
    Number3[11][12] = 4'hF;
    Number3[12][12] = 4'hF;
    Number3[13][12] = 4'hF;
    Number3[14][12] = 4'hF;
    Number3[15][12] = 4'hF;
    Number3[16][12] = 4'hF;
    Number3[17][12] = 4'hC;
    Number3[18][12] = 4'hC;
    Number3[19][12] = 4'hC;
    Number3[20][12] = 4'hC;
    Number3[21][12] = 4'hC;
    Number3[22][12] = 4'hF;
    Number3[23][12] = 4'hF;
    Number3[0][13] = 4'hF;
    Number3[1][13] = 4'hF;
    Number3[2][13] = 4'hF;
    Number3[3][13] = 4'hF;
    Number3[4][13] = 4'hF;
    Number3[5][13] = 4'hF;
    Number3[6][13] = 4'hF;
    Number3[7][13] = 4'hC;
    Number3[8][13] = 4'hC;
    Number3[9][13] = 4'hC;
    Number3[10][13] = 4'hC;
    Number3[11][13] = 4'hC;
    Number3[12][13] = 4'hC;
    Number3[13][13] = 4'hC;
    Number3[14][13] = 4'hC;
    Number3[15][13] = 4'hC;
    Number3[16][13] = 4'hC;
    Number3[17][13] = 4'hF;
    Number3[18][13] = 4'hF;
    Number3[19][13] = 4'hF;
    Number3[20][13] = 4'hF;
    Number3[21][13] = 4'hF;
    Number3[22][13] = 4'hF;
    Number3[23][13] = 4'hF;
    Number3[0][14] = 4'hF;
    Number3[1][14] = 4'hF;
    Number3[2][14] = 4'hF;
    Number3[3][14] = 4'hF;
    Number3[4][14] = 4'hF;
    Number3[5][14] = 4'hF;
    Number3[6][14] = 4'hF;
    Number3[7][14] = 4'hC;
    Number3[8][14] = 4'hC;
    Number3[9][14] = 4'hC;
    Number3[10][14] = 4'hC;
    Number3[11][14] = 4'hC;
    Number3[12][14] = 4'hC;
    Number3[13][14] = 4'hC;
    Number3[14][14] = 4'hC;
    Number3[15][14] = 4'hC;
    Number3[16][14] = 4'hC;
    Number3[17][14] = 4'hF;
    Number3[18][14] = 4'hF;
    Number3[19][14] = 4'hF;
    Number3[20][14] = 4'hF;
    Number3[21][14] = 4'hF;
    Number3[22][14] = 4'hF;
    Number3[23][14] = 4'hF;
    Number3[0][15] = 4'hF;
    Number3[1][15] = 4'hF;
    Number3[2][15] = 4'hF;
    Number3[3][15] = 4'hF;
    Number3[4][15] = 4'hF;
    Number3[5][15] = 4'hF;
    Number3[6][15] = 4'hF;
    Number3[7][15] = 4'hC;
    Number3[8][15] = 4'hC;
    Number3[9][15] = 4'hC;
    Number3[10][15] = 4'hC;
    Number3[11][15] = 4'hC;
    Number3[12][15] = 4'hC;
    Number3[13][15] = 4'hC;
    Number3[14][15] = 4'hC;
    Number3[15][15] = 4'hC;
    Number3[16][15] = 4'hC;
    Number3[17][15] = 4'hF;
    Number3[18][15] = 4'hF;
    Number3[19][15] = 4'hF;
    Number3[20][15] = 4'hF;
    Number3[21][15] = 4'hF;
    Number3[22][15] = 4'hF;
    Number3[23][15] = 4'hF;
    Number3[0][16] = 4'hF;
    Number3[1][16] = 4'hF;
    Number3[2][16] = 4'hF;
    Number3[3][16] = 4'hF;
    Number3[4][16] = 4'hF;
    Number3[5][16] = 4'hF;
    Number3[6][16] = 4'hF;
    Number3[7][16] = 4'hC;
    Number3[8][16] = 4'hC;
    Number3[9][16] = 4'hC;
    Number3[10][16] = 4'hC;
    Number3[11][16] = 4'hC;
    Number3[12][16] = 4'hC;
    Number3[13][16] = 4'hC;
    Number3[14][16] = 4'hC;
    Number3[15][16] = 4'hC;
    Number3[16][16] = 4'hC;
    Number3[17][16] = 4'hF;
    Number3[18][16] = 4'hF;
    Number3[19][16] = 4'hF;
    Number3[20][16] = 4'hF;
    Number3[21][16] = 4'hF;
    Number3[22][16] = 4'hF;
    Number3[23][16] = 4'hF;
    Number3[0][17] = 4'hF;
    Number3[1][17] = 4'hF;
    Number3[2][17] = 4'hF;
    Number3[3][17] = 4'hF;
    Number3[4][17] = 4'hF;
    Number3[5][17] = 4'hF;
    Number3[6][17] = 4'hF;
    Number3[7][17] = 4'hC;
    Number3[8][17] = 4'hC;
    Number3[9][17] = 4'hC;
    Number3[10][17] = 4'hC;
    Number3[11][17] = 4'hC;
    Number3[12][17] = 4'hC;
    Number3[13][17] = 4'hC;
    Number3[14][17] = 4'hC;
    Number3[15][17] = 4'hC;
    Number3[16][17] = 4'hC;
    Number3[17][17] = 4'hF;
    Number3[18][17] = 4'hF;
    Number3[19][17] = 4'hF;
    Number3[20][17] = 4'hF;
    Number3[21][17] = 4'hF;
    Number3[22][17] = 4'hF;
    Number3[23][17] = 4'hF;
    Number3[0][18] = 4'hF;
    Number3[1][18] = 4'hF;
    Number3[2][18] = 4'hF;
    Number3[3][18] = 4'hF;
    Number3[4][18] = 4'hF;
    Number3[5][18] = 4'hF;
    Number3[6][18] = 4'hF;
    Number3[7][18] = 4'hF;
    Number3[8][18] = 4'hF;
    Number3[9][18] = 4'hF;
    Number3[10][18] = 4'hF;
    Number3[11][18] = 4'hF;
    Number3[12][18] = 4'hF;
    Number3[13][18] = 4'hF;
    Number3[14][18] = 4'hF;
    Number3[15][18] = 4'hF;
    Number3[16][18] = 4'hF;
    Number3[17][18] = 4'hC;
    Number3[18][18] = 4'hC;
    Number3[19][18] = 4'hC;
    Number3[20][18] = 4'hC;
    Number3[21][18] = 4'hC;
    Number3[22][18] = 4'hF;
    Number3[23][18] = 4'hF;
    Number3[0][19] = 4'hF;
    Number3[1][19] = 4'hF;
    Number3[2][19] = 4'hF;
    Number3[3][19] = 4'hF;
    Number3[4][19] = 4'hF;
    Number3[5][19] = 4'hF;
    Number3[6][19] = 4'hF;
    Number3[7][19] = 4'hF;
    Number3[8][19] = 4'hF;
    Number3[9][19] = 4'hF;
    Number3[10][19] = 4'hF;
    Number3[11][19] = 4'hF;
    Number3[12][19] = 4'hF;
    Number3[13][19] = 4'hF;
    Number3[14][19] = 4'hF;
    Number3[15][19] = 4'hF;
    Number3[16][19] = 4'hF;
    Number3[17][19] = 4'hC;
    Number3[18][19] = 4'hC;
    Number3[19][19] = 4'hC;
    Number3[20][19] = 4'hC;
    Number3[21][19] = 4'hC;
    Number3[22][19] = 4'hF;
    Number3[23][19] = 4'hF;
    Number3[0][20] = 4'hF;
    Number3[1][20] = 4'hF;
    Number3[2][20] = 4'hF;
    Number3[3][20] = 4'hF;
    Number3[4][20] = 4'hF;
    Number3[5][20] = 4'hF;
    Number3[6][20] = 4'hF;
    Number3[7][20] = 4'hF;
    Number3[8][20] = 4'hF;
    Number3[9][20] = 4'hF;
    Number3[10][20] = 4'hF;
    Number3[11][20] = 4'hF;
    Number3[12][20] = 4'hF;
    Number3[13][20] = 4'hF;
    Number3[14][20] = 4'hF;
    Number3[15][20] = 4'hF;
    Number3[16][20] = 4'hF;
    Number3[17][20] = 4'hC;
    Number3[18][20] = 4'hC;
    Number3[19][20] = 4'hC;
    Number3[20][20] = 4'hC;
    Number3[21][20] = 4'hC;
    Number3[22][20] = 4'hF;
    Number3[23][20] = 4'hF;
    Number3[0][21] = 4'hF;
    Number3[1][21] = 4'hF;
    Number3[2][21] = 4'hF;
    Number3[3][21] = 4'hF;
    Number3[4][21] = 4'hF;
    Number3[5][21] = 4'hF;
    Number3[6][21] = 4'hF;
    Number3[7][21] = 4'hF;
    Number3[8][21] = 4'hF;
    Number3[9][21] = 4'hF;
    Number3[10][21] = 4'hF;
    Number3[11][21] = 4'hF;
    Number3[12][21] = 4'hF;
    Number3[13][21] = 4'hF;
    Number3[14][21] = 4'hF;
    Number3[15][21] = 4'hF;
    Number3[16][21] = 4'hF;
    Number3[17][21] = 4'hC;
    Number3[18][21] = 4'hC;
    Number3[19][21] = 4'hC;
    Number3[20][21] = 4'hC;
    Number3[21][21] = 4'hC;
    Number3[22][21] = 4'hF;
    Number3[23][21] = 4'hF;
    Number3[0][22] = 4'hF;
    Number3[1][22] = 4'hF;
    Number3[2][22] = 4'hF;
    Number3[3][22] = 4'hF;
    Number3[4][22] = 4'hF;
    Number3[5][22] = 4'hF;
    Number3[6][22] = 4'hF;
    Number3[7][22] = 4'hF;
    Number3[8][22] = 4'hF;
    Number3[9][22] = 4'hF;
    Number3[10][22] = 4'hF;
    Number3[11][22] = 4'hF;
    Number3[12][22] = 4'hF;
    Number3[13][22] = 4'hF;
    Number3[14][22] = 4'hF;
    Number3[15][22] = 4'hF;
    Number3[16][22] = 4'hF;
    Number3[17][22] = 4'hC;
    Number3[18][22] = 4'hC;
    Number3[19][22] = 4'hC;
    Number3[20][22] = 4'hC;
    Number3[21][22] = 4'hC;
    Number3[22][22] = 4'hF;
    Number3[23][22] = 4'hF;
    Number3[0][23] = 4'hF;
    Number3[1][23] = 4'hF;
    Number3[2][23] = 4'hC;
    Number3[3][23] = 4'hC;
    Number3[4][23] = 4'hC;
    Number3[5][23] = 4'hC;
    Number3[6][23] = 4'hC;
    Number3[7][23] = 4'hC;
    Number3[8][23] = 4'hC;
    Number3[9][23] = 4'hC;
    Number3[10][23] = 4'hC;
    Number3[11][23] = 4'hC;
    Number3[12][23] = 4'hC;
    Number3[13][23] = 4'hC;
    Number3[14][23] = 4'hC;
    Number3[15][23] = 4'hC;
    Number3[16][23] = 4'hC;
    Number3[17][23] = 4'hF;
    Number3[18][23] = 4'hF;
    Number3[19][23] = 4'hF;
    Number3[20][23] = 4'hF;
    Number3[21][23] = 4'hF;
    Number3[22][23] = 4'hF;
    Number3[23][23] = 4'hF;
    Number3[0][24] = 4'hF;
    Number3[1][24] = 4'hF;
    Number3[2][24] = 4'hC;
    Number3[3][24] = 4'hC;
    Number3[4][24] = 4'hC;
    Number3[5][24] = 4'hC;
    Number3[6][24] = 4'hC;
    Number3[7][24] = 4'hC;
    Number3[8][24] = 4'hC;
    Number3[9][24] = 4'hC;
    Number3[10][24] = 4'hC;
    Number3[11][24] = 4'hC;
    Number3[12][24] = 4'hC;
    Number3[13][24] = 4'hC;
    Number3[14][24] = 4'hC;
    Number3[15][24] = 4'hC;
    Number3[16][24] = 4'hC;
    Number3[17][24] = 4'hF;
    Number3[18][24] = 4'hF;
    Number3[19][24] = 4'hF;
    Number3[20][24] = 4'hF;
    Number3[21][24] = 4'hF;
    Number3[22][24] = 4'hF;
    Number3[23][24] = 4'hF;
    Number3[0][25] = 4'hF;
    Number3[1][25] = 4'hF;
    Number3[2][25] = 4'hC;
    Number3[3][25] = 4'hC;
    Number3[4][25] = 4'hC;
    Number3[5][25] = 4'hC;
    Number3[6][25] = 4'hC;
    Number3[7][25] = 4'hC;
    Number3[8][25] = 4'hC;
    Number3[9][25] = 4'hC;
    Number3[10][25] = 4'hC;
    Number3[11][25] = 4'hC;
    Number3[12][25] = 4'hC;
    Number3[13][25] = 4'hC;
    Number3[14][25] = 4'hC;
    Number3[15][25] = 4'hC;
    Number3[16][25] = 4'hC;
    Number3[17][25] = 4'hF;
    Number3[18][25] = 4'hF;
    Number3[19][25] = 4'hF;
    Number3[20][25] = 4'hF;
    Number3[21][25] = 4'hF;
    Number3[22][25] = 4'hF;
    Number3[23][25] = 4'hF;
    Number3[0][26] = 4'hF;
    Number3[1][26] = 4'hF;
    Number3[2][26] = 4'hC;
    Number3[3][26] = 4'hC;
    Number3[4][26] = 4'hC;
    Number3[5][26] = 4'hC;
    Number3[6][26] = 4'hC;
    Number3[7][26] = 4'hC;
    Number3[8][26] = 4'hC;
    Number3[9][26] = 4'hC;
    Number3[10][26] = 4'hC;
    Number3[11][26] = 4'hC;
    Number3[12][26] = 4'hC;
    Number3[13][26] = 4'hC;
    Number3[14][26] = 4'hC;
    Number3[15][26] = 4'hC;
    Number3[16][26] = 4'hC;
    Number3[17][26] = 4'hF;
    Number3[18][26] = 4'hF;
    Number3[19][26] = 4'hF;
    Number3[20][26] = 4'hF;
    Number3[21][26] = 4'hF;
    Number3[22][26] = 4'hF;
    Number3[23][26] = 4'hF;
    Number3[0][27] = 4'hF;
    Number3[1][27] = 4'hF;
    Number3[2][27] = 4'hC;
    Number3[3][27] = 4'hC;
    Number3[4][27] = 4'hC;
    Number3[5][27] = 4'hC;
    Number3[6][27] = 4'hC;
    Number3[7][27] = 4'hC;
    Number3[8][27] = 4'hC;
    Number3[9][27] = 4'hC;
    Number3[10][27] = 4'hC;
    Number3[11][27] = 4'hC;
    Number3[12][27] = 4'hC;
    Number3[13][27] = 4'hC;
    Number3[14][27] = 4'hC;
    Number3[15][27] = 4'hC;
    Number3[16][27] = 4'hC;
    Number3[17][27] = 4'hF;
    Number3[18][27] = 4'hF;
    Number3[19][27] = 4'hF;
    Number3[20][27] = 4'hF;
    Number3[21][27] = 4'hF;
    Number3[22][27] = 4'hF;
    Number3[23][27] = 4'hF;
    Number3[0][28] = 4'hF;
    Number3[1][28] = 4'hF;
    Number3[2][28] = 4'hF;
    Number3[3][28] = 4'hF;
    Number3[4][28] = 4'hF;
    Number3[5][28] = 4'hF;
    Number3[6][28] = 4'hF;
    Number3[7][28] = 4'hF;
    Number3[8][28] = 4'hF;
    Number3[9][28] = 4'hF;
    Number3[10][28] = 4'hF;
    Number3[11][28] = 4'hF;
    Number3[12][28] = 4'hF;
    Number3[13][28] = 4'hF;
    Number3[14][28] = 4'hF;
    Number3[15][28] = 4'hF;
    Number3[16][28] = 4'hF;
    Number3[17][28] = 4'hF;
    Number3[18][28] = 4'hF;
    Number3[19][28] = 4'hF;
    Number3[20][28] = 4'hF;
    Number3[21][28] = 4'hF;
    Number3[22][28] = 4'hF;
    Number3[23][28] = 4'hF;
    Number3[0][29] = 4'hF;
    Number3[1][29] = 4'hF;
    Number3[2][29] = 4'hF;
    Number3[3][29] = 4'hF;
    Number3[4][29] = 4'hF;
    Number3[5][29] = 4'hF;
    Number3[6][29] = 4'hF;
    Number3[7][29] = 4'hF;
    Number3[8][29] = 4'hF;
    Number3[9][29] = 4'hF;
    Number3[10][29] = 4'hF;
    Number3[11][29] = 4'hF;
    Number3[12][29] = 4'hF;
    Number3[13][29] = 4'hF;
    Number3[14][29] = 4'hF;
    Number3[15][29] = 4'hF;
    Number3[16][29] = 4'hF;
    Number3[17][29] = 4'hF;
    Number3[18][29] = 4'hF;
    Number3[19][29] = 4'hF;
    Number3[20][29] = 4'hF;
    Number3[21][29] = 4'hF;
    Number3[22][29] = 4'hF;
    Number3[23][29] = 4'hF;
 
//Number 4
    Number4[0][0] = 4'hF;
    Number4[1][0] = 4'hF;
    Number4[2][0] = 4'hF;
    Number4[3][0] = 4'hF;
    Number4[4][0] = 4'hF;
    Number4[5][0] = 4'hF;
    Number4[6][0] = 4'hF;
    Number4[7][0] = 4'hF;
    Number4[8][0] = 4'hF;
    Number4[9][0] = 4'hF;
    Number4[10][0] = 4'hF;
    Number4[11][0] = 4'hF;
    Number4[12][0] = 4'hF;
    Number4[13][0] = 4'hF;
    Number4[14][0] = 4'hF;
    Number4[15][0] = 4'hF;
    Number4[16][0] = 4'hF;
    Number4[17][0] = 4'hF;
    Number4[18][0] = 4'hF;
    Number4[19][0] = 4'hF;
    Number4[20][0] = 4'hF;
    Number4[21][0] = 4'hF;
    Number4[22][0] = 4'hF;
    Number4[23][0] = 4'hF;
    Number4[0][1] = 4'hF;
    Number4[1][1] = 4'hF;
    Number4[2][1] = 4'hF;
    Number4[3][1] = 4'hF;
    Number4[4][1] = 4'hF;
    Number4[5][1] = 4'hF;
    Number4[6][1] = 4'hF;
    Number4[7][1] = 4'hF;
    Number4[8][1] = 4'hF;
    Number4[9][1] = 4'hF;
    Number4[10][1] = 4'hF;
    Number4[11][1] = 4'hF;
    Number4[12][1] = 4'hF;
    Number4[13][1] = 4'hF;
    Number4[14][1] = 4'hF;
    Number4[15][1] = 4'hF;
    Number4[16][1] = 4'hF;
    Number4[17][1] = 4'hF;
    Number4[18][1] = 4'hF;
    Number4[19][1] = 4'hF;
    Number4[20][1] = 4'hF;
    Number4[21][1] = 4'hF;
    Number4[22][1] = 4'hF;
    Number4[23][1] = 4'hF;
    Number4[0][2] = 4'hF;
    Number4[1][2] = 4'hF;
    Number4[2][2] = 4'hF;
    Number4[3][2] = 4'hF;
    Number4[4][2] = 4'hF;
    Number4[5][2] = 4'hF;
    Number4[6][2] = 4'hF;
    Number4[7][2] = 4'hF;
    Number4[8][2] = 4'hF;
    Number4[9][2] = 4'hF;
    Number4[10][2] = 4'hF;
    Number4[11][2] = 4'hF;
    Number4[12][2] = 4'hF;
    Number4[13][2] = 4'hF;
    Number4[14][2] = 4'hF;
    Number4[15][2] = 4'hF;
    Number4[16][2] = 4'hF;
    Number4[17][2] = 4'hF;
    Number4[18][2] = 4'hF;
    Number4[19][2] = 4'hF;
    Number4[20][2] = 4'hF;
    Number4[21][2] = 4'hF;
    Number4[22][2] = 4'hF;
    Number4[23][2] = 4'hF;
    Number4[0][3] = 4'hF;
    Number4[1][3] = 4'hF;
    Number4[2][3] = 4'hF;
    Number4[3][3] = 4'hF;
    Number4[4][3] = 4'hF;
    Number4[5][3] = 4'hF;
    Number4[6][3] = 4'hF;
    Number4[7][3] = 4'hF;
    Number4[8][3] = 4'hF;
    Number4[9][3] = 4'hF;
    Number4[10][3] = 4'hF;
    Number4[11][3] = 4'hF;
    Number4[12][3] = 4'hC;
    Number4[13][3] = 4'hC;
    Number4[14][3] = 4'hC;
    Number4[15][3] = 4'hC;
    Number4[16][3] = 4'hC;
    Number4[17][3] = 4'hF;
    Number4[18][3] = 4'hF;
    Number4[19][3] = 4'hF;
    Number4[20][3] = 4'hF;
    Number4[21][3] = 4'hF;
    Number4[22][3] = 4'hF;
    Number4[23][3] = 4'hF;
    Number4[0][4] = 4'hF;
    Number4[1][4] = 4'hF;
    Number4[2][4] = 4'hF;
    Number4[3][4] = 4'hF;
    Number4[4][4] = 4'hF;
    Number4[5][4] = 4'hF;
    Number4[6][4] = 4'hF;
    Number4[7][4] = 4'hF;
    Number4[8][4] = 4'hF;
    Number4[9][4] = 4'hF;
    Number4[10][4] = 4'hF;
    Number4[11][4] = 4'hF;
    Number4[12][4] = 4'hC;
    Number4[13][4] = 4'hC;
    Number4[14][4] = 4'hC;
    Number4[15][4] = 4'hC;
    Number4[16][4] = 4'hC;
    Number4[17][4] = 4'hF;
    Number4[18][4] = 4'hF;
    Number4[19][4] = 4'hF;
    Number4[20][4] = 4'hF;
    Number4[21][4] = 4'hF;
    Number4[22][4] = 4'hF;
    Number4[23][4] = 4'hF;
    Number4[0][5] = 4'hF;
    Number4[1][5] = 4'hF;
    Number4[2][5] = 4'hF;
    Number4[3][5] = 4'hF;
    Number4[4][5] = 4'hF;
    Number4[5][5] = 4'hF;
    Number4[6][5] = 4'hF;
    Number4[7][5] = 4'hF;
    Number4[8][5] = 4'hF;
    Number4[9][5] = 4'hF;
    Number4[10][5] = 4'hF;
    Number4[11][5] = 4'hF;
    Number4[12][5] = 4'hC;
    Number4[13][5] = 4'hC;
    Number4[14][5] = 4'hC;
    Number4[15][5] = 4'hC;
    Number4[16][5] = 4'hC;
    Number4[17][5] = 4'hF;
    Number4[18][5] = 4'hF;
    Number4[19][5] = 4'hF;
    Number4[20][5] = 4'hF;
    Number4[21][5] = 4'hF;
    Number4[22][5] = 4'hF;
    Number4[23][5] = 4'hF;
    Number4[0][6] = 4'hF;
    Number4[1][6] = 4'hF;
    Number4[2][6] = 4'hF;
    Number4[3][6] = 4'hF;
    Number4[4][6] = 4'hF;
    Number4[5][6] = 4'hF;
    Number4[6][6] = 4'hF;
    Number4[7][6] = 4'hF;
    Number4[8][6] = 4'hF;
    Number4[9][6] = 4'hF;
    Number4[10][6] = 4'hF;
    Number4[11][6] = 4'hF;
    Number4[12][6] = 4'hC;
    Number4[13][6] = 4'hC;
    Number4[14][6] = 4'hC;
    Number4[15][6] = 4'hC;
    Number4[16][6] = 4'hC;
    Number4[17][6] = 4'hF;
    Number4[18][6] = 4'hF;
    Number4[19][6] = 4'hF;
    Number4[20][6] = 4'hF;
    Number4[21][6] = 4'hF;
    Number4[22][6] = 4'hF;
    Number4[23][6] = 4'hF;
    Number4[0][7] = 4'hF;
    Number4[1][7] = 4'hF;
    Number4[2][7] = 4'hF;
    Number4[3][7] = 4'hF;
    Number4[4][7] = 4'hF;
    Number4[5][7] = 4'hF;
    Number4[6][7] = 4'hF;
    Number4[7][7] = 4'hF;
    Number4[8][7] = 4'hF;
    Number4[9][7] = 4'hF;
    Number4[10][7] = 4'hF;
    Number4[11][7] = 4'hF;
    Number4[12][7] = 4'hC;
    Number4[13][7] = 4'hC;
    Number4[14][7] = 4'hC;
    Number4[15][7] = 4'hC;
    Number4[16][7] = 4'hC;
    Number4[17][7] = 4'hF;
    Number4[18][7] = 4'hF;
    Number4[19][7] = 4'hF;
    Number4[20][7] = 4'hF;
    Number4[21][7] = 4'hF;
    Number4[22][7] = 4'hF;
    Number4[23][7] = 4'hF;
    Number4[0][8] = 4'hF;
    Number4[1][8] = 4'hF;
    Number4[2][8] = 4'hF;
    Number4[3][8] = 4'hF;
    Number4[4][8] = 4'hF;
    Number4[5][8] = 4'hF;
    Number4[6][8] = 4'hF;
    Number4[7][8] = 4'hC;
    Number4[8][8] = 4'hC;
    Number4[9][8] = 4'hC;
    Number4[10][8] = 4'hC;
    Number4[11][8] = 4'hC;
    Number4[12][8] = 4'hC;
    Number4[13][8] = 4'hC;
    Number4[14][8] = 4'hC;
    Number4[15][8] = 4'hC;
    Number4[16][8] = 4'hC;
    Number4[17][8] = 4'hF;
    Number4[18][8] = 4'hF;
    Number4[19][8] = 4'hF;
    Number4[20][8] = 4'hF;
    Number4[21][8] = 4'hF;
    Number4[22][8] = 4'hF;
    Number4[23][8] = 4'hF;
    Number4[0][9] = 4'hF;
    Number4[1][9] = 4'hF;
    Number4[2][9] = 4'hF;
    Number4[3][9] = 4'hF;
    Number4[4][9] = 4'hF;
    Number4[5][9] = 4'hF;
    Number4[6][9] = 4'hF;
    Number4[7][9] = 4'hC;
    Number4[8][9] = 4'hC;
    Number4[9][9] = 4'hC;
    Number4[10][9] = 4'hC;
    Number4[11][9] = 4'hC;
    Number4[12][9] = 4'hC;
    Number4[13][9] = 4'hC;
    Number4[14][9] = 4'hC;
    Number4[15][9] = 4'hC;
    Number4[16][9] = 4'hC;
    Number4[17][9] = 4'hF;
    Number4[18][9] = 4'hF;
    Number4[19][9] = 4'hF;
    Number4[20][9] = 4'hF;
    Number4[21][9] = 4'hF;
    Number4[22][9] = 4'hF;
    Number4[23][9] = 4'hF;
    Number4[0][10] = 4'hF;
    Number4[1][10] = 4'hF;
    Number4[2][10] = 4'hF;
    Number4[3][10] = 4'hF;
    Number4[4][10] = 4'hF;
    Number4[5][10] = 4'hF;
    Number4[6][10] = 4'hF;
    Number4[7][10] = 4'hC;
    Number4[8][10] = 4'hC;
    Number4[9][10] = 4'hC;
    Number4[10][10] = 4'hC;
    Number4[11][10] = 4'hC;
    Number4[12][10] = 4'hC;
    Number4[13][10] = 4'hC;
    Number4[14][10] = 4'hC;
    Number4[15][10] = 4'hC;
    Number4[16][10] = 4'hC;
    Number4[17][10] = 4'hF;
    Number4[18][10] = 4'hF;
    Number4[19][10] = 4'hF;
    Number4[20][10] = 4'hF;
    Number4[21][10] = 4'hF;
    Number4[22][10] = 4'hF;
    Number4[23][10] = 4'hF;
    Number4[0][11] = 4'hF;
    Number4[1][11] = 4'hF;
    Number4[2][11] = 4'hF;
    Number4[3][11] = 4'hF;
    Number4[4][11] = 4'hF;
    Number4[5][11] = 4'hF;
    Number4[6][11] = 4'hF;
    Number4[7][11] = 4'hC;
    Number4[8][11] = 4'hC;
    Number4[9][11] = 4'hC;
    Number4[10][11] = 4'hC;
    Number4[11][11] = 4'hC;
    Number4[12][11] = 4'hC;
    Number4[13][11] = 4'hC;
    Number4[14][11] = 4'hC;
    Number4[15][11] = 4'hC;
    Number4[16][11] = 4'hC;
    Number4[17][11] = 4'hF;
    Number4[18][11] = 4'hF;
    Number4[19][11] = 4'hF;
    Number4[20][11] = 4'hF;
    Number4[21][11] = 4'hF;
    Number4[22][11] = 4'hF;
    Number4[23][11] = 4'hF;
    Number4[0][12] = 4'hF;
    Number4[1][12] = 4'hF;
    Number4[2][12] = 4'hF;
    Number4[3][12] = 4'hF;
    Number4[4][12] = 4'hF;
    Number4[5][12] = 4'hF;
    Number4[6][12] = 4'hF;
    Number4[7][12] = 4'hC;
    Number4[8][12] = 4'hC;
    Number4[9][12] = 4'hC;
    Number4[10][12] = 4'hC;
    Number4[11][12] = 4'hC;
    Number4[12][12] = 4'hC;
    Number4[13][12] = 4'hC;
    Number4[14][12] = 4'hC;
    Number4[15][12] = 4'hC;
    Number4[16][12] = 4'hC;
    Number4[17][12] = 4'hF;
    Number4[18][12] = 4'hF;
    Number4[19][12] = 4'hF;
    Number4[20][12] = 4'hF;
    Number4[21][12] = 4'hF;
    Number4[22][12] = 4'hF;
    Number4[23][12] = 4'hF;
    Number4[0][13] = 4'hF;
    Number4[1][13] = 4'hF;
    Number4[2][13] = 4'hC;
    Number4[3][13] = 4'hC;
    Number4[4][13] = 4'hC;
    Number4[5][13] = 4'hC;
    Number4[6][13] = 4'hC;
    Number4[7][13] = 4'hF;
    Number4[8][13] = 4'hF;
    Number4[9][13] = 4'hF;
    Number4[10][13] = 4'hF;
    Number4[11][13] = 4'hF;
    Number4[12][13] = 4'hC;
    Number4[13][13] = 4'hC;
    Number4[14][13] = 4'hC;
    Number4[15][13] = 4'hC;
    Number4[16][13] = 4'hC;
    Number4[17][13] = 4'hF;
    Number4[18][13] = 4'hF;
    Number4[19][13] = 4'hF;
    Number4[20][13] = 4'hF;
    Number4[21][13] = 4'hF;
    Number4[22][13] = 4'hF;
    Number4[23][13] = 4'hF;
    Number4[0][14] = 4'hF;
    Number4[1][14] = 4'hF;
    Number4[2][14] = 4'hC;
    Number4[3][14] = 4'hC;
    Number4[4][14] = 4'hC;
    Number4[5][14] = 4'hC;
    Number4[6][14] = 4'hC;
    Number4[7][14] = 4'hF;
    Number4[8][14] = 4'hF;
    Number4[9][14] = 4'hF;
    Number4[10][14] = 4'hF;
    Number4[11][14] = 4'hF;
    Number4[12][14] = 4'hC;
    Number4[13][14] = 4'hC;
    Number4[14][14] = 4'hC;
    Number4[15][14] = 4'hC;
    Number4[16][14] = 4'hC;
    Number4[17][14] = 4'hF;
    Number4[18][14] = 4'hF;
    Number4[19][14] = 4'hF;
    Number4[20][14] = 4'hF;
    Number4[21][14] = 4'hF;
    Number4[22][14] = 4'hF;
    Number4[23][14] = 4'hF;
    Number4[0][15] = 4'hF;
    Number4[1][15] = 4'hF;
    Number4[2][15] = 4'hC;
    Number4[3][15] = 4'hC;
    Number4[4][15] = 4'hC;
    Number4[5][15] = 4'hC;
    Number4[6][15] = 4'hC;
    Number4[7][15] = 4'hF;
    Number4[8][15] = 4'hF;
    Number4[9][15] = 4'hF;
    Number4[10][15] = 4'hF;
    Number4[11][15] = 4'hF;
    Number4[12][15] = 4'hC;
    Number4[13][15] = 4'hC;
    Number4[14][15] = 4'hC;
    Number4[15][15] = 4'hC;
    Number4[16][15] = 4'hC;
    Number4[17][15] = 4'hF;
    Number4[18][15] = 4'hF;
    Number4[19][15] = 4'hF;
    Number4[20][15] = 4'hF;
    Number4[21][15] = 4'hF;
    Number4[22][15] = 4'hF;
    Number4[23][15] = 4'hF;
    Number4[0][16] = 4'hF;
    Number4[1][16] = 4'hF;
    Number4[2][16] = 4'hC;
    Number4[3][16] = 4'hC;
    Number4[4][16] = 4'hC;
    Number4[5][16] = 4'hC;
    Number4[6][16] = 4'hC;
    Number4[7][16] = 4'hF;
    Number4[8][16] = 4'hF;
    Number4[9][16] = 4'hF;
    Number4[10][16] = 4'hF;
    Number4[11][16] = 4'hF;
    Number4[12][16] = 4'hC;
    Number4[13][16] = 4'hC;
    Number4[14][16] = 4'hC;
    Number4[15][16] = 4'hC;
    Number4[16][16] = 4'hC;
    Number4[17][16] = 4'hF;
    Number4[18][16] = 4'hF;
    Number4[19][16] = 4'hF;
    Number4[20][16] = 4'hF;
    Number4[21][16] = 4'hF;
    Number4[22][16] = 4'hF;
    Number4[23][16] = 4'hF;
    Number4[0][17] = 4'hF;
    Number4[1][17] = 4'hF;
    Number4[2][17] = 4'hC;
    Number4[3][17] = 4'hC;
    Number4[4][17] = 4'hC;
    Number4[5][17] = 4'hC;
    Number4[6][17] = 4'hC;
    Number4[7][17] = 4'hF;
    Number4[8][17] = 4'hF;
    Number4[9][17] = 4'hF;
    Number4[10][17] = 4'hF;
    Number4[11][17] = 4'hF;
    Number4[12][17] = 4'hC;
    Number4[13][17] = 4'hC;
    Number4[14][17] = 4'hC;
    Number4[15][17] = 4'hC;
    Number4[16][17] = 4'hC;
    Number4[17][17] = 4'hF;
    Number4[18][17] = 4'hF;
    Number4[19][17] = 4'hF;
    Number4[20][17] = 4'hF;
    Number4[21][17] = 4'hF;
    Number4[22][17] = 4'hF;
    Number4[23][17] = 4'hF;
    Number4[0][18] = 4'hF;
    Number4[1][18] = 4'hF;
    Number4[2][18] = 4'hC;
    Number4[3][18] = 4'hC;
    Number4[4][18] = 4'hC;
    Number4[5][18] = 4'hC;
    Number4[6][18] = 4'hC;
    Number4[7][18] = 4'hC;
    Number4[8][18] = 4'hC;
    Number4[9][18] = 4'hC;
    Number4[10][18] = 4'hC;
    Number4[11][18] = 4'hC;
    Number4[12][18] = 4'hC;
    Number4[13][18] = 4'hC;
    Number4[14][18] = 4'hC;
    Number4[15][18] = 4'hC;
    Number4[16][18] = 4'hC;
    Number4[17][18] = 4'hC;
    Number4[18][18] = 4'hC;
    Number4[19][18] = 4'hC;
    Number4[20][18] = 4'hC;
    Number4[21][18] = 4'hC;
    Number4[22][18] = 4'hF;
    Number4[23][18] = 4'hF;
    Number4[0][19] = 4'hF;
    Number4[1][19] = 4'hF;
    Number4[2][19] = 4'hC;
    Number4[3][19] = 4'hC;
    Number4[4][19] = 4'hC;
    Number4[5][19] = 4'hC;
    Number4[6][19] = 4'hC;
    Number4[7][19] = 4'hC;
    Number4[8][19] = 4'hC;
    Number4[9][19] = 4'hC;
    Number4[10][19] = 4'hC;
    Number4[11][19] = 4'hC;
    Number4[12][19] = 4'hC;
    Number4[13][19] = 4'hC;
    Number4[14][19] = 4'hC;
    Number4[15][19] = 4'hC;
    Number4[16][19] = 4'hC;
    Number4[17][19] = 4'hC;
    Number4[18][19] = 4'hC;
    Number4[19][19] = 4'hC;
    Number4[20][19] = 4'hC;
    Number4[21][19] = 4'hC;
    Number4[22][19] = 4'hF;
    Number4[23][19] = 4'hF;
    Number4[0][20] = 4'hF;
    Number4[1][20] = 4'hF;
    Number4[2][20] = 4'hC;
    Number4[3][20] = 4'hC;
    Number4[4][20] = 4'hC;
    Number4[5][20] = 4'hC;
    Number4[6][20] = 4'hC;
    Number4[7][20] = 4'hC;
    Number4[8][20] = 4'hC;
    Number4[9][20] = 4'hC;
    Number4[10][20] = 4'hC;
    Number4[11][20] = 4'hC;
    Number4[12][20] = 4'hC;
    Number4[13][20] = 4'hC;
    Number4[14][20] = 4'hC;
    Number4[15][20] = 4'hC;
    Number4[16][20] = 4'hC;
    Number4[17][20] = 4'hC;
    Number4[18][20] = 4'hC;
    Number4[19][20] = 4'hC;
    Number4[20][20] = 4'hC;
    Number4[21][20] = 4'hC;
    Number4[22][20] = 4'hF;
    Number4[23][20] = 4'hF;
    Number4[0][21] = 4'hF;
    Number4[1][21] = 4'hF;
    Number4[2][21] = 4'hC;
    Number4[3][21] = 4'hC;
    Number4[4][21] = 4'hC;
    Number4[5][21] = 4'hC;
    Number4[6][21] = 4'hC;
    Number4[7][21] = 4'hC;
    Number4[8][21] = 4'hC;
    Number4[9][21] = 4'hC;
    Number4[10][21] = 4'hC;
    Number4[11][21] = 4'hC;
    Number4[12][21] = 4'hC;
    Number4[13][21] = 4'hC;
    Number4[14][21] = 4'hC;
    Number4[15][21] = 4'hC;
    Number4[16][21] = 4'hC;
    Number4[17][21] = 4'hC;
    Number4[18][21] = 4'hC;
    Number4[19][21] = 4'hC;
    Number4[20][21] = 4'hC;
    Number4[21][21] = 4'hC;
    Number4[22][21] = 4'hF;
    Number4[23][21] = 4'hF;
    Number4[0][22] = 4'hF;
    Number4[1][22] = 4'hF;
    Number4[2][22] = 4'hC;
    Number4[3][22] = 4'hC;
    Number4[4][22] = 4'hC;
    Number4[5][22] = 4'hC;
    Number4[6][22] = 4'hC;
    Number4[7][22] = 4'hC;
    Number4[8][22] = 4'hC;
    Number4[9][22] = 4'hC;
    Number4[10][22] = 4'hC;
    Number4[11][22] = 4'hC;
    Number4[12][22] = 4'hC;
    Number4[13][22] = 4'hC;
    Number4[14][22] = 4'hC;
    Number4[15][22] = 4'hC;
    Number4[16][22] = 4'hC;
    Number4[17][22] = 4'hC;
    Number4[18][22] = 4'hC;
    Number4[19][22] = 4'hC;
    Number4[20][22] = 4'hC;
    Number4[21][22] = 4'hC;
    Number4[22][22] = 4'hF;
    Number4[23][22] = 4'hF;
    Number4[0][23] = 4'hF;
    Number4[1][23] = 4'hF;
    Number4[2][23] = 4'hF;
    Number4[3][23] = 4'hF;
    Number4[4][23] = 4'hF;
    Number4[5][23] = 4'hF;
    Number4[6][23] = 4'hF;
    Number4[7][23] = 4'hF;
    Number4[8][23] = 4'hF;
    Number4[9][23] = 4'hF;
    Number4[10][23] = 4'hF;
    Number4[11][23] = 4'hF;
    Number4[12][23] = 4'hC;
    Number4[13][23] = 4'hC;
    Number4[14][23] = 4'hC;
    Number4[15][23] = 4'hC;
    Number4[16][23] = 4'hC;
    Number4[17][23] = 4'hF;
    Number4[18][23] = 4'hF;
    Number4[19][23] = 4'hF;
    Number4[20][23] = 4'hF;
    Number4[21][23] = 4'hF;
    Number4[22][23] = 4'hF;
    Number4[23][23] = 4'hF;
    Number4[0][24] = 4'hF;
    Number4[1][24] = 4'hF;
    Number4[2][24] = 4'hF;
    Number4[3][24] = 4'hF;
    Number4[4][24] = 4'hF;
    Number4[5][24] = 4'hF;
    Number4[6][24] = 4'hF;
    Number4[7][24] = 4'hF;
    Number4[8][24] = 4'hF;
    Number4[9][24] = 4'hF;
    Number4[10][24] = 4'hF;
    Number4[11][24] = 4'hF;
    Number4[12][24] = 4'hC;
    Number4[13][24] = 4'hC;
    Number4[14][24] = 4'hC;
    Number4[15][24] = 4'hC;
    Number4[16][24] = 4'hC;
    Number4[17][24] = 4'hF;
    Number4[18][24] = 4'hF;
    Number4[19][24] = 4'hF;
    Number4[20][24] = 4'hF;
    Number4[21][24] = 4'hF;
    Number4[22][24] = 4'hF;
    Number4[23][24] = 4'hF;
    Number4[0][25] = 4'hF;
    Number4[1][25] = 4'hF;
    Number4[2][25] = 4'hF;
    Number4[3][25] = 4'hF;
    Number4[4][25] = 4'hF;
    Number4[5][25] = 4'hF;
    Number4[6][25] = 4'hF;
    Number4[7][25] = 4'hF;
    Number4[8][25] = 4'hF;
    Number4[9][25] = 4'hF;
    Number4[10][25] = 4'hF;
    Number4[11][25] = 4'hF;
    Number4[12][25] = 4'hC;
    Number4[13][25] = 4'hC;
    Number4[14][25] = 4'hC;
    Number4[15][25] = 4'hC;
    Number4[16][25] = 4'hC;
    Number4[17][25] = 4'hF;
    Number4[18][25] = 4'hF;
    Number4[19][25] = 4'hF;
    Number4[20][25] = 4'hF;
    Number4[21][25] = 4'hF;
    Number4[22][25] = 4'hF;
    Number4[23][25] = 4'hF;
    Number4[0][26] = 4'hF;
    Number4[1][26] = 4'hF;
    Number4[2][26] = 4'hF;
    Number4[3][26] = 4'hF;
    Number4[4][26] = 4'hF;
    Number4[5][26] = 4'hF;
    Number4[6][26] = 4'hF;
    Number4[7][26] = 4'hF;
    Number4[8][26] = 4'hF;
    Number4[9][26] = 4'hF;
    Number4[10][26] = 4'hF;
    Number4[11][26] = 4'hF;
    Number4[12][26] = 4'hC;
    Number4[13][26] = 4'hC;
    Number4[14][26] = 4'hC;
    Number4[15][26] = 4'hC;
    Number4[16][26] = 4'hC;
    Number4[17][26] = 4'hF;
    Number4[18][26] = 4'hF;
    Number4[19][26] = 4'hF;
    Number4[20][26] = 4'hF;
    Number4[21][26] = 4'hF;
    Number4[22][26] = 4'hF;
    Number4[23][26] = 4'hF;
    Number4[0][27] = 4'hF;
    Number4[1][27] = 4'hF;
    Number4[2][27] = 4'hF;
    Number4[3][27] = 4'hF;
    Number4[4][27] = 4'hF;
    Number4[5][27] = 4'hF;
    Number4[6][27] = 4'hF;
    Number4[7][27] = 4'hF;
    Number4[8][27] = 4'hF;
    Number4[9][27] = 4'hF;
    Number4[10][27] = 4'hF;
    Number4[11][27] = 4'hF;
    Number4[12][27] = 4'hC;
    Number4[13][27] = 4'hC;
    Number4[14][27] = 4'hC;
    Number4[15][27] = 4'hC;
    Number4[16][27] = 4'hC;
    Number4[17][27] = 4'hF;
    Number4[18][27] = 4'hF;
    Number4[19][27] = 4'hF;
    Number4[20][27] = 4'hF;
    Number4[21][27] = 4'hF;
    Number4[22][27] = 4'hF;
    Number4[23][27] = 4'hF;
    Number4[0][28] = 4'hF;
    Number4[1][28] = 4'hF;
    Number4[2][28] = 4'hF;
    Number4[3][28] = 4'hF;
    Number4[4][28] = 4'hF;
    Number4[5][28] = 4'hF;
    Number4[6][28] = 4'hF;
    Number4[7][28] = 4'hF;
    Number4[8][28] = 4'hF;
    Number4[9][28] = 4'hF;
    Number4[10][28] = 4'hF;
    Number4[11][28] = 4'hF;
    Number4[12][28] = 4'hF;
    Number4[13][28] = 4'hF;
    Number4[14][28] = 4'hF;
    Number4[15][28] = 4'hF;
    Number4[16][28] = 4'hF;
    Number4[17][28] = 4'hF;
    Number4[18][28] = 4'hF;
    Number4[19][28] = 4'hF;
    Number4[20][28] = 4'hF;
    Number4[21][28] = 4'hF;
    Number4[22][28] = 4'hF;
    Number4[23][28] = 4'hF;
    Number4[0][29] = 4'hF;
    Number4[1][29] = 4'hF;
    Number4[2][29] = 4'hF;
    Number4[3][29] = 4'hF;
    Number4[4][29] = 4'hF;
    Number4[5][29] = 4'hF;
    Number4[6][29] = 4'hF;
    Number4[7][29] = 4'hF;
    Number4[8][29] = 4'hF;
    Number4[9][29] = 4'hF;
    Number4[10][29] = 4'hF;
    Number4[11][29] = 4'hF;
    Number4[12][29] = 4'hF;
    Number4[13][29] = 4'hF;
    Number4[14][29] = 4'hF;
    Number4[15][29] = 4'hF;
    Number4[16][29] = 4'hF;
    Number4[17][29] = 4'hF;
    Number4[18][29] = 4'hF;
    Number4[19][29] = 4'hF;
    Number4[20][29] = 4'hF;
    Number4[21][29] = 4'hF;
    Number4[22][29] = 4'hF;
    Number4[23][29] = 4'hF;
 
//Number 5
    Number5[0][0] = 4'hF;
    Number5[1][0] = 4'hF;
    Number5[2][0] = 4'hF;
    Number5[3][0] = 4'hF;
    Number5[4][0] = 4'hF;
    Number5[5][0] = 4'hF;
    Number5[6][0] = 4'hF;
    Number5[7][0] = 4'hF;
    Number5[8][0] = 4'hF;
    Number5[9][0] = 4'hF;
    Number5[10][0] = 4'hF;
    Number5[11][0] = 4'hF;
    Number5[12][0] = 4'hF;
    Number5[13][0] = 4'hF;
    Number5[14][0] = 4'hF;
    Number5[15][0] = 4'hF;
    Number5[16][0] = 4'hF;
    Number5[17][0] = 4'hF;
    Number5[18][0] = 4'hF;
    Number5[19][0] = 4'hF;
    Number5[20][0] = 4'hF;
    Number5[21][0] = 4'hF;
    Number5[22][0] = 4'hF;
    Number5[23][0] = 4'hF;
    Number5[0][1] = 4'hF;
    Number5[1][1] = 4'hF;
    Number5[2][1] = 4'hF;
    Number5[3][1] = 4'hF;
    Number5[4][1] = 4'hF;
    Number5[5][1] = 4'hF;
    Number5[6][1] = 4'hF;
    Number5[7][1] = 4'hF;
    Number5[8][1] = 4'hF;
    Number5[9][1] = 4'hF;
    Number5[10][1] = 4'hF;
    Number5[11][1] = 4'hF;
    Number5[12][1] = 4'hF;
    Number5[13][1] = 4'hF;
    Number5[14][1] = 4'hF;
    Number5[15][1] = 4'hF;
    Number5[16][1] = 4'hF;
    Number5[17][1] = 4'hF;
    Number5[18][1] = 4'hF;
    Number5[19][1] = 4'hF;
    Number5[20][1] = 4'hF;
    Number5[21][1] = 4'hF;
    Number5[22][1] = 4'hF;
    Number5[23][1] = 4'hF;
    Number5[0][2] = 4'hF;
    Number5[1][2] = 4'hF;
    Number5[2][2] = 4'hF;
    Number5[3][2] = 4'hF;
    Number5[4][2] = 4'hF;
    Number5[5][2] = 4'hF;
    Number5[6][2] = 4'hF;
    Number5[7][2] = 4'hF;
    Number5[8][2] = 4'hF;
    Number5[9][2] = 4'hF;
    Number5[10][2] = 4'hF;
    Number5[11][2] = 4'hF;
    Number5[12][2] = 4'hF;
    Number5[13][2] = 4'hF;
    Number5[14][2] = 4'hF;
    Number5[15][2] = 4'hF;
    Number5[16][2] = 4'hF;
    Number5[17][2] = 4'hF;
    Number5[18][2] = 4'hF;
    Number5[19][2] = 4'hF;
    Number5[20][2] = 4'hF;
    Number5[21][2] = 4'hF;
    Number5[22][2] = 4'hF;
    Number5[23][2] = 4'hF;
    Number5[0][3] = 4'hF;
    Number5[1][3] = 4'hF;
    Number5[2][3] = 4'hC;
    Number5[3][3] = 4'hC;
    Number5[4][3] = 4'hC;
    Number5[5][3] = 4'hC;
    Number5[6][3] = 4'hC;
    Number5[7][3] = 4'hC;
    Number5[8][3] = 4'hC;
    Number5[9][3] = 4'hC;
    Number5[10][3] = 4'hC;
    Number5[11][3] = 4'hC;
    Number5[12][3] = 4'hC;
    Number5[13][3] = 4'hC;
    Number5[14][3] = 4'hC;
    Number5[15][3] = 4'hC;
    Number5[16][3] = 4'hC;
    Number5[17][3] = 4'hC;
    Number5[18][3] = 4'hC;
    Number5[19][3] = 4'hC;
    Number5[20][3] = 4'hC;
    Number5[21][3] = 4'hC;
    Number5[22][3] = 4'hF;
    Number5[23][3] = 4'hF;
    Number5[0][4] = 4'hF;
    Number5[1][4] = 4'hF;
    Number5[2][4] = 4'hC;
    Number5[3][4] = 4'hC;
    Number5[4][4] = 4'hC;
    Number5[5][4] = 4'hC;
    Number5[6][4] = 4'hC;
    Number5[7][4] = 4'hC;
    Number5[8][4] = 4'hC;
    Number5[9][4] = 4'hC;
    Number5[10][4] = 4'hC;
    Number5[11][4] = 4'hC;
    Number5[12][4] = 4'hC;
    Number5[13][4] = 4'hC;
    Number5[14][4] = 4'hC;
    Number5[15][4] = 4'hC;
    Number5[16][4] = 4'hC;
    Number5[17][4] = 4'hC;
    Number5[18][4] = 4'hC;
    Number5[19][4] = 4'hC;
    Number5[20][4] = 4'hC;
    Number5[21][4] = 4'hC;
    Number5[22][4] = 4'hF;
    Number5[23][4] = 4'hF;
    Number5[0][5] = 4'hF;
    Number5[1][5] = 4'hF;
    Number5[2][5] = 4'hC;
    Number5[3][5] = 4'hC;
    Number5[4][5] = 4'hC;
    Number5[5][5] = 4'hC;
    Number5[6][5] = 4'hC;
    Number5[7][5] = 4'hC;
    Number5[8][5] = 4'hC;
    Number5[9][5] = 4'hC;
    Number5[10][5] = 4'hC;
    Number5[11][5] = 4'hC;
    Number5[12][5] = 4'hC;
    Number5[13][5] = 4'hC;
    Number5[14][5] = 4'hC;
    Number5[15][5] = 4'hC;
    Number5[16][5] = 4'hC;
    Number5[17][5] = 4'hC;
    Number5[18][5] = 4'hC;
    Number5[19][5] = 4'hC;
    Number5[20][5] = 4'hC;
    Number5[21][5] = 4'hC;
    Number5[22][5] = 4'hF;
    Number5[23][5] = 4'hF;
    Number5[0][6] = 4'hF;
    Number5[1][6] = 4'hF;
    Number5[2][6] = 4'hC;
    Number5[3][6] = 4'hC;
    Number5[4][6] = 4'hC;
    Number5[5][6] = 4'hC;
    Number5[6][6] = 4'hC;
    Number5[7][6] = 4'hC;
    Number5[8][6] = 4'hC;
    Number5[9][6] = 4'hC;
    Number5[10][6] = 4'hC;
    Number5[11][6] = 4'hC;
    Number5[12][6] = 4'hC;
    Number5[13][6] = 4'hC;
    Number5[14][6] = 4'hC;
    Number5[15][6] = 4'hC;
    Number5[16][6] = 4'hC;
    Number5[17][6] = 4'hC;
    Number5[18][6] = 4'hC;
    Number5[19][6] = 4'hC;
    Number5[20][6] = 4'hC;
    Number5[21][6] = 4'hC;
    Number5[22][6] = 4'hF;
    Number5[23][6] = 4'hF;
    Number5[0][7] = 4'hF;
    Number5[1][7] = 4'hF;
    Number5[2][7] = 4'hC;
    Number5[3][7] = 4'hC;
    Number5[4][7] = 4'hC;
    Number5[5][7] = 4'hC;
    Number5[6][7] = 4'hC;
    Number5[7][7] = 4'hC;
    Number5[8][7] = 4'hC;
    Number5[9][7] = 4'hC;
    Number5[10][7] = 4'hC;
    Number5[11][7] = 4'hC;
    Number5[12][7] = 4'hC;
    Number5[13][7] = 4'hC;
    Number5[14][7] = 4'hC;
    Number5[15][7] = 4'hC;
    Number5[16][7] = 4'hC;
    Number5[17][7] = 4'hC;
    Number5[18][7] = 4'hC;
    Number5[19][7] = 4'hC;
    Number5[20][7] = 4'hC;
    Number5[21][7] = 4'hC;
    Number5[22][7] = 4'hF;
    Number5[23][7] = 4'hF;
    Number5[0][8] = 4'hF;
    Number5[1][8] = 4'hF;
    Number5[2][8] = 4'hC;
    Number5[3][8] = 4'hC;
    Number5[4][8] = 4'hC;
    Number5[5][8] = 4'hC;
    Number5[6][8] = 4'hC;
    Number5[7][8] = 4'hF;
    Number5[8][8] = 4'hF;
    Number5[9][8] = 4'hF;
    Number5[10][8] = 4'hF;
    Number5[11][8] = 4'hF;
    Number5[12][8] = 4'hF;
    Number5[13][8] = 4'hF;
    Number5[14][8] = 4'hF;
    Number5[15][8] = 4'hF;
    Number5[16][8] = 4'hF;
    Number5[17][8] = 4'hF;
    Number5[18][8] = 4'hF;
    Number5[19][8] = 4'hF;
    Number5[20][8] = 4'hF;
    Number5[21][8] = 4'hF;
    Number5[22][8] = 4'hF;
    Number5[23][8] = 4'hF;
    Number5[0][9] = 4'hF;
    Number5[1][9] = 4'hF;
    Number5[2][9] = 4'hC;
    Number5[3][9] = 4'hC;
    Number5[4][9] = 4'hC;
    Number5[5][9] = 4'hC;
    Number5[6][9] = 4'hC;
    Number5[7][9] = 4'hF;
    Number5[8][9] = 4'hF;
    Number5[9][9] = 4'hF;
    Number5[10][9] = 4'hF;
    Number5[11][9] = 4'hF;
    Number5[12][9] = 4'hF;
    Number5[13][9] = 4'hF;
    Number5[14][9] = 4'hF;
    Number5[15][9] = 4'hF;
    Number5[16][9] = 4'hF;
    Number5[17][9] = 4'hF;
    Number5[18][9] = 4'hF;
    Number5[19][9] = 4'hF;
    Number5[20][9] = 4'hF;
    Number5[21][9] = 4'hF;
    Number5[22][9] = 4'hF;
    Number5[23][9] = 4'hF;
    Number5[0][10] = 4'hF;
    Number5[1][10] = 4'hF;
    Number5[2][10] = 4'hC;
    Number5[3][10] = 4'hC;
    Number5[4][10] = 4'hC;
    Number5[5][10] = 4'hC;
    Number5[6][10] = 4'hC;
    Number5[7][10] = 4'hF;
    Number5[8][10] = 4'hF;
    Number5[9][10] = 4'hF;
    Number5[10][10] = 4'hF;
    Number5[11][10] = 4'hF;
    Number5[12][10] = 4'hF;
    Number5[13][10] = 4'hF;
    Number5[14][10] = 4'hF;
    Number5[15][10] = 4'hF;
    Number5[16][10] = 4'hF;
    Number5[17][10] = 4'hF;
    Number5[18][10] = 4'hF;
    Number5[19][10] = 4'hF;
    Number5[20][10] = 4'hF;
    Number5[21][10] = 4'hF;
    Number5[22][10] = 4'hF;
    Number5[23][10] = 4'hF;
    Number5[0][11] = 4'hF;
    Number5[1][11] = 4'hF;
    Number5[2][11] = 4'hC;
    Number5[3][11] = 4'hC;
    Number5[4][11] = 4'hC;
    Number5[5][11] = 4'hC;
    Number5[6][11] = 4'hC;
    Number5[7][11] = 4'hF;
    Number5[8][11] = 4'hF;
    Number5[9][11] = 4'hF;
    Number5[10][11] = 4'hF;
    Number5[11][11] = 4'hF;
    Number5[12][11] = 4'hF;
    Number5[13][11] = 4'hF;
    Number5[14][11] = 4'hF;
    Number5[15][11] = 4'hF;
    Number5[16][11] = 4'hF;
    Number5[17][11] = 4'hF;
    Number5[18][11] = 4'hF;
    Number5[19][11] = 4'hF;
    Number5[20][11] = 4'hF;
    Number5[21][11] = 4'hF;
    Number5[22][11] = 4'hF;
    Number5[23][11] = 4'hF;
    Number5[0][12] = 4'hF;
    Number5[1][12] = 4'hF;
    Number5[2][12] = 4'hC;
    Number5[3][12] = 4'hC;
    Number5[4][12] = 4'hC;
    Number5[5][12] = 4'hC;
    Number5[6][12] = 4'hC;
    Number5[7][12] = 4'hF;
    Number5[8][12] = 4'hF;
    Number5[9][12] = 4'hF;
    Number5[10][12] = 4'hF;
    Number5[11][12] = 4'hF;
    Number5[12][12] = 4'hF;
    Number5[13][12] = 4'hF;
    Number5[14][12] = 4'hF;
    Number5[15][12] = 4'hF;
    Number5[16][12] = 4'hF;
    Number5[17][12] = 4'hF;
    Number5[18][12] = 4'hF;
    Number5[19][12] = 4'hF;
    Number5[20][12] = 4'hF;
    Number5[21][12] = 4'hF;
    Number5[22][12] = 4'hF;
    Number5[23][12] = 4'hF;
    Number5[0][13] = 4'hF;
    Number5[1][13] = 4'hF;
    Number5[2][13] = 4'hC;
    Number5[3][13] = 4'hC;
    Number5[4][13] = 4'hC;
    Number5[5][13] = 4'hC;
    Number5[6][13] = 4'hC;
    Number5[7][13] = 4'hC;
    Number5[8][13] = 4'hC;
    Number5[9][13] = 4'hC;
    Number5[10][13] = 4'hC;
    Number5[11][13] = 4'hC;
    Number5[12][13] = 4'hC;
    Number5[13][13] = 4'hC;
    Number5[14][13] = 4'hC;
    Number5[15][13] = 4'hC;
    Number5[16][13] = 4'hC;
    Number5[17][13] = 4'hF;
    Number5[18][13] = 4'hF;
    Number5[19][13] = 4'hF;
    Number5[20][13] = 4'hF;
    Number5[21][13] = 4'hF;
    Number5[22][13] = 4'hF;
    Number5[23][13] = 4'hF;
    Number5[0][14] = 4'hF;
    Number5[1][14] = 4'hF;
    Number5[2][14] = 4'hC;
    Number5[3][14] = 4'hC;
    Number5[4][14] = 4'hC;
    Number5[5][14] = 4'hC;
    Number5[6][14] = 4'hC;
    Number5[7][14] = 4'hC;
    Number5[8][14] = 4'hC;
    Number5[9][14] = 4'hC;
    Number5[10][14] = 4'hC;
    Number5[11][14] = 4'hC;
    Number5[12][14] = 4'hC;
    Number5[13][14] = 4'hC;
    Number5[14][14] = 4'hC;
    Number5[15][14] = 4'hC;
    Number5[16][14] = 4'hC;
    Number5[17][14] = 4'hF;
    Number5[18][14] = 4'hF;
    Number5[19][14] = 4'hF;
    Number5[20][14] = 4'hF;
    Number5[21][14] = 4'hF;
    Number5[22][14] = 4'hF;
    Number5[23][14] = 4'hF;
    Number5[0][15] = 4'hF;
    Number5[1][15] = 4'hF;
    Number5[2][15] = 4'hC;
    Number5[3][15] = 4'hC;
    Number5[4][15] = 4'hC;
    Number5[5][15] = 4'hC;
    Number5[6][15] = 4'hC;
    Number5[7][15] = 4'hC;
    Number5[8][15] = 4'hC;
    Number5[9][15] = 4'hC;
    Number5[10][15] = 4'hC;
    Number5[11][15] = 4'hC;
    Number5[12][15] = 4'hC;
    Number5[13][15] = 4'hC;
    Number5[14][15] = 4'hC;
    Number5[15][15] = 4'hC;
    Number5[16][15] = 4'hC;
    Number5[17][15] = 4'hF;
    Number5[18][15] = 4'hF;
    Number5[19][15] = 4'hF;
    Number5[20][15] = 4'hF;
    Number5[21][15] = 4'hF;
    Number5[22][15] = 4'hF;
    Number5[23][15] = 4'hF;
    Number5[0][16] = 4'hF;
    Number5[1][16] = 4'hF;
    Number5[2][16] = 4'hC;
    Number5[3][16] = 4'hC;
    Number5[4][16] = 4'hC;
    Number5[5][16] = 4'hC;
    Number5[6][16] = 4'hC;
    Number5[7][16] = 4'hC;
    Number5[8][16] = 4'hC;
    Number5[9][16] = 4'hC;
    Number5[10][16] = 4'hC;
    Number5[11][16] = 4'hC;
    Number5[12][16] = 4'hC;
    Number5[13][16] = 4'hC;
    Number5[14][16] = 4'hC;
    Number5[15][16] = 4'hC;
    Number5[16][16] = 4'hC;
    Number5[17][16] = 4'hF;
    Number5[18][16] = 4'hF;
    Number5[19][16] = 4'hF;
    Number5[20][16] = 4'hF;
    Number5[21][16] = 4'hF;
    Number5[22][16] = 4'hF;
    Number5[23][16] = 4'hF;
    Number5[0][17] = 4'hF;
    Number5[1][17] = 4'hF;
    Number5[2][17] = 4'hC;
    Number5[3][17] = 4'hC;
    Number5[4][17] = 4'hC;
    Number5[5][17] = 4'hC;
    Number5[6][17] = 4'hC;
    Number5[7][17] = 4'hC;
    Number5[8][17] = 4'hC;
    Number5[9][17] = 4'hC;
    Number5[10][17] = 4'hC;
    Number5[11][17] = 4'hC;
    Number5[12][17] = 4'hC;
    Number5[13][17] = 4'hC;
    Number5[14][17] = 4'hC;
    Number5[15][17] = 4'hC;
    Number5[16][17] = 4'hC;
    Number5[17][17] = 4'hF;
    Number5[18][17] = 4'hF;
    Number5[19][17] = 4'hF;
    Number5[20][17] = 4'hF;
    Number5[21][17] = 4'hF;
    Number5[22][17] = 4'hF;
    Number5[23][17] = 4'hF;
    Number5[0][18] = 4'hF;
    Number5[1][18] = 4'hF;
    Number5[2][18] = 4'hF;
    Number5[3][18] = 4'hF;
    Number5[4][18] = 4'hF;
    Number5[5][18] = 4'hF;
    Number5[6][18] = 4'hF;
    Number5[7][18] = 4'hF;
    Number5[8][18] = 4'hF;
    Number5[9][18] = 4'hF;
    Number5[10][18] = 4'hF;
    Number5[11][18] = 4'hF;
    Number5[12][18] = 4'hF;
    Number5[13][18] = 4'hF;
    Number5[14][18] = 4'hF;
    Number5[15][18] = 4'hF;
    Number5[16][18] = 4'hF;
    Number5[17][18] = 4'hC;
    Number5[18][18] = 4'hC;
    Number5[19][18] = 4'hC;
    Number5[20][18] = 4'hC;
    Number5[21][18] = 4'hC;
    Number5[22][18] = 4'hF;
    Number5[23][18] = 4'hF;
    Number5[0][19] = 4'hF;
    Number5[1][19] = 4'hF;
    Number5[2][19] = 4'hF;
    Number5[3][19] = 4'hF;
    Number5[4][19] = 4'hF;
    Number5[5][19] = 4'hF;
    Number5[6][19] = 4'hF;
    Number5[7][19] = 4'hF;
    Number5[8][19] = 4'hF;
    Number5[9][19] = 4'hF;
    Number5[10][19] = 4'hF;
    Number5[11][19] = 4'hF;
    Number5[12][19] = 4'hF;
    Number5[13][19] = 4'hF;
    Number5[14][19] = 4'hF;
    Number5[15][19] = 4'hF;
    Number5[16][19] = 4'hF;
    Number5[17][19] = 4'hC;
    Number5[18][19] = 4'hC;
    Number5[19][19] = 4'hC;
    Number5[20][19] = 4'hC;
    Number5[21][19] = 4'hC;
    Number5[22][19] = 4'hF;
    Number5[23][19] = 4'hF;
    Number5[0][20] = 4'hF;
    Number5[1][20] = 4'hF;
    Number5[2][20] = 4'hF;
    Number5[3][20] = 4'hF;
    Number5[4][20] = 4'hF;
    Number5[5][20] = 4'hF;
    Number5[6][20] = 4'hF;
    Number5[7][20] = 4'hF;
    Number5[8][20] = 4'hF;
    Number5[9][20] = 4'hF;
    Number5[10][20] = 4'hF;
    Number5[11][20] = 4'hF;
    Number5[12][20] = 4'hF;
    Number5[13][20] = 4'hF;
    Number5[14][20] = 4'hF;
    Number5[15][20] = 4'hF;
    Number5[16][20] = 4'hF;
    Number5[17][20] = 4'hC;
    Number5[18][20] = 4'hC;
    Number5[19][20] = 4'hC;
    Number5[20][20] = 4'hC;
    Number5[21][20] = 4'hC;
    Number5[22][20] = 4'hF;
    Number5[23][20] = 4'hF;
    Number5[0][21] = 4'hF;
    Number5[1][21] = 4'hF;
    Number5[2][21] = 4'hF;
    Number5[3][21] = 4'hF;
    Number5[4][21] = 4'hF;
    Number5[5][21] = 4'hF;
    Number5[6][21] = 4'hF;
    Number5[7][21] = 4'hF;
    Number5[8][21] = 4'hF;
    Number5[9][21] = 4'hF;
    Number5[10][21] = 4'hF;
    Number5[11][21] = 4'hF;
    Number5[12][21] = 4'hF;
    Number5[13][21] = 4'hF;
    Number5[14][21] = 4'hF;
    Number5[15][21] = 4'hF;
    Number5[16][21] = 4'hF;
    Number5[17][21] = 4'hC;
    Number5[18][21] = 4'hC;
    Number5[19][21] = 4'hC;
    Number5[20][21] = 4'hC;
    Number5[21][21] = 4'hC;
    Number5[22][21] = 4'hF;
    Number5[23][21] = 4'hF;
    Number5[0][22] = 4'hF;
    Number5[1][22] = 4'hF;
    Number5[2][22] = 4'hF;
    Number5[3][22] = 4'hF;
    Number5[4][22] = 4'hF;
    Number5[5][22] = 4'hF;
    Number5[6][22] = 4'hF;
    Number5[7][22] = 4'hF;
    Number5[8][22] = 4'hF;
    Number5[9][22] = 4'hF;
    Number5[10][22] = 4'hF;
    Number5[11][22] = 4'hF;
    Number5[12][22] = 4'hF;
    Number5[13][22] = 4'hF;
    Number5[14][22] = 4'hF;
    Number5[15][22] = 4'hF;
    Number5[16][22] = 4'hF;
    Number5[17][22] = 4'hC;
    Number5[18][22] = 4'hC;
    Number5[19][22] = 4'hC;
    Number5[20][22] = 4'hC;
    Number5[21][22] = 4'hC;
    Number5[22][22] = 4'hF;
    Number5[23][22] = 4'hF;
    Number5[0][23] = 4'hF;
    Number5[1][23] = 4'hF;
    Number5[2][23] = 4'hC;
    Number5[3][23] = 4'hC;
    Number5[4][23] = 4'hC;
    Number5[5][23] = 4'hC;
    Number5[6][23] = 4'hC;
    Number5[7][23] = 4'hC;
    Number5[8][23] = 4'hC;
    Number5[9][23] = 4'hC;
    Number5[10][23] = 4'hC;
    Number5[11][23] = 4'hC;
    Number5[12][23] = 4'hC;
    Number5[13][23] = 4'hC;
    Number5[14][23] = 4'hC;
    Number5[15][23] = 4'hC;
    Number5[16][23] = 4'hC;
    Number5[17][23] = 4'hF;
    Number5[18][23] = 4'hF;
    Number5[19][23] = 4'hF;
    Number5[20][23] = 4'hF;
    Number5[21][23] = 4'hF;
    Number5[22][23] = 4'hF;
    Number5[23][23] = 4'hF;
    Number5[0][24] = 4'hF;
    Number5[1][24] = 4'hF;
    Number5[2][24] = 4'hC;
    Number5[3][24] = 4'hC;
    Number5[4][24] = 4'hC;
    Number5[5][24] = 4'hC;
    Number5[6][24] = 4'hC;
    Number5[7][24] = 4'hC;
    Number5[8][24] = 4'hC;
    Number5[9][24] = 4'hC;
    Number5[10][24] = 4'hC;
    Number5[11][24] = 4'hC;
    Number5[12][24] = 4'hC;
    Number5[13][24] = 4'hC;
    Number5[14][24] = 4'hC;
    Number5[15][24] = 4'hC;
    Number5[16][24] = 4'hC;
    Number5[17][24] = 4'hF;
    Number5[18][24] = 4'hF;
    Number5[19][24] = 4'hF;
    Number5[20][24] = 4'hF;
    Number5[21][24] = 4'hF;
    Number5[22][24] = 4'hF;
    Number5[23][24] = 4'hF;
    Number5[0][25] = 4'hF;
    Number5[1][25] = 4'hF;
    Number5[2][25] = 4'hC;
    Number5[3][25] = 4'hC;
    Number5[4][25] = 4'hC;
    Number5[5][25] = 4'hC;
    Number5[6][25] = 4'hC;
    Number5[7][25] = 4'hC;
    Number5[8][25] = 4'hC;
    Number5[9][25] = 4'hC;
    Number5[10][25] = 4'hC;
    Number5[11][25] = 4'hC;
    Number5[12][25] = 4'hC;
    Number5[13][25] = 4'hC;
    Number5[14][25] = 4'hC;
    Number5[15][25] = 4'hC;
    Number5[16][25] = 4'hC;
    Number5[17][25] = 4'hF;
    Number5[18][25] = 4'hF;
    Number5[19][25] = 4'hF;
    Number5[20][25] = 4'hF;
    Number5[21][25] = 4'hF;
    Number5[22][25] = 4'hF;
    Number5[23][25] = 4'hF;
    Number5[0][26] = 4'hF;
    Number5[1][26] = 4'hF;
    Number5[2][26] = 4'hC;
    Number5[3][26] = 4'hC;
    Number5[4][26] = 4'hC;
    Number5[5][26] = 4'hC;
    Number5[6][26] = 4'hC;
    Number5[7][26] = 4'hC;
    Number5[8][26] = 4'hC;
    Number5[9][26] = 4'hC;
    Number5[10][26] = 4'hC;
    Number5[11][26] = 4'hC;
    Number5[12][26] = 4'hC;
    Number5[13][26] = 4'hC;
    Number5[14][26] = 4'hC;
    Number5[15][26] = 4'hC;
    Number5[16][26] = 4'hC;
    Number5[17][26] = 4'hF;
    Number5[18][26] = 4'hF;
    Number5[19][26] = 4'hF;
    Number5[20][26] = 4'hF;
    Number5[21][26] = 4'hF;
    Number5[22][26] = 4'hF;
    Number5[23][26] = 4'hF;
    Number5[0][27] = 4'hF;
    Number5[1][27] = 4'hF;
    Number5[2][27] = 4'hC;
    Number5[3][27] = 4'hC;
    Number5[4][27] = 4'hC;
    Number5[5][27] = 4'hC;
    Number5[6][27] = 4'hC;
    Number5[7][27] = 4'hC;
    Number5[8][27] = 4'hC;
    Number5[9][27] = 4'hC;
    Number5[10][27] = 4'hC;
    Number5[11][27] = 4'hC;
    Number5[12][27] = 4'hC;
    Number5[13][27] = 4'hC;
    Number5[14][27] = 4'hC;
    Number5[15][27] = 4'hC;
    Number5[16][27] = 4'hC;
    Number5[17][27] = 4'hF;
    Number5[18][27] = 4'hF;
    Number5[19][27] = 4'hF;
    Number5[20][27] = 4'hF;
    Number5[21][27] = 4'hF;
    Number5[22][27] = 4'hF;
    Number5[23][27] = 4'hF;
    Number5[0][28] = 4'hF;
    Number5[1][28] = 4'hF;
    Number5[2][28] = 4'hF;
    Number5[3][28] = 4'hF;
    Number5[4][28] = 4'hF;
    Number5[5][28] = 4'hF;
    Number5[6][28] = 4'hF;
    Number5[7][28] = 4'hF;
    Number5[8][28] = 4'hF;
    Number5[9][28] = 4'hF;
    Number5[10][28] = 4'hF;
    Number5[11][28] = 4'hF;
    Number5[12][28] = 4'hF;
    Number5[13][28] = 4'hF;
    Number5[14][28] = 4'hF;
    Number5[15][28] = 4'hF;
    Number5[16][28] = 4'hF;
    Number5[17][28] = 4'hF;
    Number5[18][28] = 4'hF;
    Number5[19][28] = 4'hF;
    Number5[20][28] = 4'hF;
    Number5[21][28] = 4'hF;
    Number5[22][28] = 4'hF;
    Number5[23][28] = 4'hF;
    Number5[0][29] = 4'hF;
    Number5[1][29] = 4'hF;
    Number5[2][29] = 4'hF;
    Number5[3][29] = 4'hF;
    Number5[4][29] = 4'hF;
    Number5[5][29] = 4'hF;
    Number5[6][29] = 4'hF;
    Number5[7][29] = 4'hF;
    Number5[8][29] = 4'hF;
    Number5[9][29] = 4'hF;
    Number5[10][29] = 4'hF;
    Number5[11][29] = 4'hF;
    Number5[12][29] = 4'hF;
    Number5[13][29] = 4'hF;
    Number5[14][29] = 4'hF;
    Number5[15][29] = 4'hF;
    Number5[16][29] = 4'hF;
    Number5[17][29] = 4'hF;
    Number5[18][29] = 4'hF;
    Number5[19][29] = 4'hF;
    Number5[20][29] = 4'hF;
    Number5[21][29] = 4'hF;
    Number5[22][29] = 4'hF;
    Number5[23][29] = 4'hF;
 
//Number 6
    Number6[0][0] = 4'hF;
    Number6[1][0] = 4'hF;
    Number6[2][0] = 4'hF;
    Number6[3][0] = 4'hF;
    Number6[4][0] = 4'hF;
    Number6[5][0] = 4'hF;
    Number6[6][0] = 4'hF;
    Number6[7][0] = 4'hF;
    Number6[8][0] = 4'hF;
    Number6[9][0] = 4'hF;
    Number6[10][0] = 4'hF;
    Number6[11][0] = 4'hF;
    Number6[12][0] = 4'hF;
    Number6[13][0] = 4'hF;
    Number6[14][0] = 4'hF;
    Number6[15][0] = 4'hF;
    Number6[16][0] = 4'hF;
    Number6[17][0] = 4'hF;
    Number6[18][0] = 4'hF;
    Number6[19][0] = 4'hF;
    Number6[20][0] = 4'hF;
    Number6[21][0] = 4'hF;
    Number6[22][0] = 4'hF;
    Number6[23][0] = 4'hF;
    Number6[0][1] = 4'hF;
    Number6[1][1] = 4'hF;
    Number6[2][1] = 4'hF;
    Number6[3][1] = 4'hF;
    Number6[4][1] = 4'hF;
    Number6[5][1] = 4'hF;
    Number6[6][1] = 4'hF;
    Number6[7][1] = 4'hF;
    Number6[8][1] = 4'hF;
    Number6[9][1] = 4'hF;
    Number6[10][1] = 4'hF;
    Number6[11][1] = 4'hF;
    Number6[12][1] = 4'hF;
    Number6[13][1] = 4'hF;
    Number6[14][1] = 4'hF;
    Number6[15][1] = 4'hF;
    Number6[16][1] = 4'hF;
    Number6[17][1] = 4'hF;
    Number6[18][1] = 4'hF;
    Number6[19][1] = 4'hF;
    Number6[20][1] = 4'hF;
    Number6[21][1] = 4'hF;
    Number6[22][1] = 4'hF;
    Number6[23][1] = 4'hF;
    Number6[0][2] = 4'hF;
    Number6[1][2] = 4'hF;
    Number6[2][2] = 4'hF;
    Number6[3][2] = 4'hF;
    Number6[4][2] = 4'hF;
    Number6[5][2] = 4'hF;
    Number6[6][2] = 4'hF;
    Number6[7][2] = 4'hF;
    Number6[8][2] = 4'hF;
    Number6[9][2] = 4'hF;
    Number6[10][2] = 4'hF;
    Number6[11][2] = 4'hF;
    Number6[12][2] = 4'hF;
    Number6[13][2] = 4'hF;
    Number6[14][2] = 4'hF;
    Number6[15][2] = 4'hF;
    Number6[16][2] = 4'hF;
    Number6[17][2] = 4'hF;
    Number6[18][2] = 4'hF;
    Number6[19][2] = 4'hF;
    Number6[20][2] = 4'hF;
    Number6[21][2] = 4'hF;
    Number6[22][2] = 4'hF;
    Number6[23][2] = 4'hF;
    Number6[0][3] = 4'hF;
    Number6[1][3] = 4'hF;
    Number6[2][3] = 4'hF;
    Number6[3][3] = 4'hF;
    Number6[4][3] = 4'hF;
    Number6[5][3] = 4'hF;
    Number6[6][3] = 4'hF;
    Number6[7][3] = 4'hC;
    Number6[8][3] = 4'hC;
    Number6[9][3] = 4'hC;
    Number6[10][3] = 4'hC;
    Number6[11][3] = 4'hC;
    Number6[12][3] = 4'hC;
    Number6[13][3] = 4'hC;
    Number6[14][3] = 4'hC;
    Number6[15][3] = 4'hC;
    Number6[16][3] = 4'hC;
    Number6[17][3] = 4'hF;
    Number6[18][3] = 4'hF;
    Number6[19][3] = 4'hF;
    Number6[20][3] = 4'hF;
    Number6[21][3] = 4'hF;
    Number6[22][3] = 4'hF;
    Number6[23][3] = 4'hF;
    Number6[0][4] = 4'hF;
    Number6[1][4] = 4'hF;
    Number6[2][4] = 4'hF;
    Number6[3][4] = 4'hF;
    Number6[4][4] = 4'hF;
    Number6[5][4] = 4'hF;
    Number6[6][4] = 4'hF;
    Number6[7][4] = 4'hC;
    Number6[8][4] = 4'hC;
    Number6[9][4] = 4'hC;
    Number6[10][4] = 4'hC;
    Number6[11][4] = 4'hC;
    Number6[12][4] = 4'hC;
    Number6[13][4] = 4'hC;
    Number6[14][4] = 4'hC;
    Number6[15][4] = 4'hC;
    Number6[16][4] = 4'hC;
    Number6[17][4] = 4'hF;
    Number6[18][4] = 4'hF;
    Number6[19][4] = 4'hF;
    Number6[20][4] = 4'hF;
    Number6[21][4] = 4'hF;
    Number6[22][4] = 4'hF;
    Number6[23][4] = 4'hF;
    Number6[0][5] = 4'hF;
    Number6[1][5] = 4'hF;
    Number6[2][5] = 4'hF;
    Number6[3][5] = 4'hF;
    Number6[4][5] = 4'hF;
    Number6[5][5] = 4'hF;
    Number6[6][5] = 4'hF;
    Number6[7][5] = 4'hC;
    Number6[8][5] = 4'hC;
    Number6[9][5] = 4'hC;
    Number6[10][5] = 4'hC;
    Number6[11][5] = 4'hC;
    Number6[12][5] = 4'hC;
    Number6[13][5] = 4'hC;
    Number6[14][5] = 4'hC;
    Number6[15][5] = 4'hC;
    Number6[16][5] = 4'hC;
    Number6[17][5] = 4'hF;
    Number6[18][5] = 4'hF;
    Number6[19][5] = 4'hF;
    Number6[20][5] = 4'hF;
    Number6[21][5] = 4'hF;
    Number6[22][5] = 4'hF;
    Number6[23][5] = 4'hF;
    Number6[0][6] = 4'hF;
    Number6[1][6] = 4'hF;
    Number6[2][6] = 4'hF;
    Number6[3][6] = 4'hF;
    Number6[4][6] = 4'hF;
    Number6[5][6] = 4'hF;
    Number6[6][6] = 4'hF;
    Number6[7][6] = 4'hC;
    Number6[8][6] = 4'hC;
    Number6[9][6] = 4'hC;
    Number6[10][6] = 4'hC;
    Number6[11][6] = 4'hC;
    Number6[12][6] = 4'hC;
    Number6[13][6] = 4'hC;
    Number6[14][6] = 4'hC;
    Number6[15][6] = 4'hC;
    Number6[16][6] = 4'hC;
    Number6[17][6] = 4'hF;
    Number6[18][6] = 4'hF;
    Number6[19][6] = 4'hF;
    Number6[20][6] = 4'hF;
    Number6[21][6] = 4'hF;
    Number6[22][6] = 4'hF;
    Number6[23][6] = 4'hF;
    Number6[0][7] = 4'hF;
    Number6[1][7] = 4'hF;
    Number6[2][7] = 4'hF;
    Number6[3][7] = 4'hF;
    Number6[4][7] = 4'hF;
    Number6[5][7] = 4'hF;
    Number6[6][7] = 4'hF;
    Number6[7][7] = 4'hC;
    Number6[8][7] = 4'hC;
    Number6[9][7] = 4'hC;
    Number6[10][7] = 4'hC;
    Number6[11][7] = 4'hC;
    Number6[12][7] = 4'hC;
    Number6[13][7] = 4'hC;
    Number6[14][7] = 4'hC;
    Number6[15][7] = 4'hC;
    Number6[16][7] = 4'hC;
    Number6[17][7] = 4'hF;
    Number6[18][7] = 4'hF;
    Number6[19][7] = 4'hF;
    Number6[20][7] = 4'hF;
    Number6[21][7] = 4'hF;
    Number6[22][7] = 4'hF;
    Number6[23][7] = 4'hF;
    Number6[0][8] = 4'hF;
    Number6[1][8] = 4'hF;
    Number6[2][8] = 4'hC;
    Number6[3][8] = 4'hC;
    Number6[4][8] = 4'hC;
    Number6[5][8] = 4'hC;
    Number6[6][8] = 4'hC;
    Number6[7][8] = 4'hF;
    Number6[8][8] = 4'hF;
    Number6[9][8] = 4'hF;
    Number6[10][8] = 4'hF;
    Number6[11][8] = 4'hF;
    Number6[12][8] = 4'hF;
    Number6[13][8] = 4'hF;
    Number6[14][8] = 4'hF;
    Number6[15][8] = 4'hF;
    Number6[16][8] = 4'hF;
    Number6[17][8] = 4'hF;
    Number6[18][8] = 4'hF;
    Number6[19][8] = 4'hF;
    Number6[20][8] = 4'hF;
    Number6[21][8] = 4'hF;
    Number6[22][8] = 4'hF;
    Number6[23][8] = 4'hF;
    Number6[0][9] = 4'hF;
    Number6[1][9] = 4'hF;
    Number6[2][9] = 4'hC;
    Number6[3][9] = 4'hC;
    Number6[4][9] = 4'hC;
    Number6[5][9] = 4'hC;
    Number6[6][9] = 4'hC;
    Number6[7][9] = 4'hF;
    Number6[8][9] = 4'hF;
    Number6[9][9] = 4'hF;
    Number6[10][9] = 4'hF;
    Number6[11][9] = 4'hF;
    Number6[12][9] = 4'hF;
    Number6[13][9] = 4'hF;
    Number6[14][9] = 4'hF;
    Number6[15][9] = 4'hF;
    Number6[16][9] = 4'hF;
    Number6[17][9] = 4'hF;
    Number6[18][9] = 4'hF;
    Number6[19][9] = 4'hF;
    Number6[20][9] = 4'hF;
    Number6[21][9] = 4'hF;
    Number6[22][9] = 4'hF;
    Number6[23][9] = 4'hF;
    Number6[0][10] = 4'hF;
    Number6[1][10] = 4'hF;
    Number6[2][10] = 4'hC;
    Number6[3][10] = 4'hC;
    Number6[4][10] = 4'hC;
    Number6[5][10] = 4'hC;
    Number6[6][10] = 4'hC;
    Number6[7][10] = 4'hF;
    Number6[8][10] = 4'hF;
    Number6[9][10] = 4'hF;
    Number6[10][10] = 4'hF;
    Number6[11][10] = 4'hF;
    Number6[12][10] = 4'hF;
    Number6[13][10] = 4'hF;
    Number6[14][10] = 4'hF;
    Number6[15][10] = 4'hF;
    Number6[16][10] = 4'hF;
    Number6[17][10] = 4'hF;
    Number6[18][10] = 4'hF;
    Number6[19][10] = 4'hF;
    Number6[20][10] = 4'hF;
    Number6[21][10] = 4'hF;
    Number6[22][10] = 4'hF;
    Number6[23][10] = 4'hF;
    Number6[0][11] = 4'hF;
    Number6[1][11] = 4'hF;
    Number6[2][11] = 4'hC;
    Number6[3][11] = 4'hC;
    Number6[4][11] = 4'hC;
    Number6[5][11] = 4'hC;
    Number6[6][11] = 4'hC;
    Number6[7][11] = 4'hF;
    Number6[8][11] = 4'hF;
    Number6[9][11] = 4'hF;
    Number6[10][11] = 4'hF;
    Number6[11][11] = 4'hF;
    Number6[12][11] = 4'hF;
    Number6[13][11] = 4'hF;
    Number6[14][11] = 4'hF;
    Number6[15][11] = 4'hF;
    Number6[16][11] = 4'hF;
    Number6[17][11] = 4'hF;
    Number6[18][11] = 4'hF;
    Number6[19][11] = 4'hF;
    Number6[20][11] = 4'hF;
    Number6[21][11] = 4'hF;
    Number6[22][11] = 4'hF;
    Number6[23][11] = 4'hF;
    Number6[0][12] = 4'hF;
    Number6[1][12] = 4'hF;
    Number6[2][12] = 4'hC;
    Number6[3][12] = 4'hC;
    Number6[4][12] = 4'hC;
    Number6[5][12] = 4'hC;
    Number6[6][12] = 4'hC;
    Number6[7][12] = 4'hF;
    Number6[8][12] = 4'hF;
    Number6[9][12] = 4'hF;
    Number6[10][12] = 4'hF;
    Number6[11][12] = 4'hF;
    Number6[12][12] = 4'hF;
    Number6[13][12] = 4'hF;
    Number6[14][12] = 4'hF;
    Number6[15][12] = 4'hF;
    Number6[16][12] = 4'hF;
    Number6[17][12] = 4'hF;
    Number6[18][12] = 4'hF;
    Number6[19][12] = 4'hF;
    Number6[20][12] = 4'hF;
    Number6[21][12] = 4'hF;
    Number6[22][12] = 4'hF;
    Number6[23][12] = 4'hF;
    Number6[0][13] = 4'hF;
    Number6[1][13] = 4'hF;
    Number6[2][13] = 4'hC;
    Number6[3][13] = 4'hC;
    Number6[4][13] = 4'hC;
    Number6[5][13] = 4'hC;
    Number6[6][13] = 4'hC;
    Number6[7][13] = 4'hC;
    Number6[8][13] = 4'hC;
    Number6[9][13] = 4'hC;
    Number6[10][13] = 4'hC;
    Number6[11][13] = 4'hC;
    Number6[12][13] = 4'hC;
    Number6[13][13] = 4'hC;
    Number6[14][13] = 4'hC;
    Number6[15][13] = 4'hC;
    Number6[16][13] = 4'hC;
    Number6[17][13] = 4'hF;
    Number6[18][13] = 4'hF;
    Number6[19][13] = 4'hF;
    Number6[20][13] = 4'hF;
    Number6[21][13] = 4'hF;
    Number6[22][13] = 4'hF;
    Number6[23][13] = 4'hF;
    Number6[0][14] = 4'hF;
    Number6[1][14] = 4'hF;
    Number6[2][14] = 4'hC;
    Number6[3][14] = 4'hC;
    Number6[4][14] = 4'hC;
    Number6[5][14] = 4'hC;
    Number6[6][14] = 4'hC;
    Number6[7][14] = 4'hC;
    Number6[8][14] = 4'hC;
    Number6[9][14] = 4'hC;
    Number6[10][14] = 4'hC;
    Number6[11][14] = 4'hC;
    Number6[12][14] = 4'hC;
    Number6[13][14] = 4'hC;
    Number6[14][14] = 4'hC;
    Number6[15][14] = 4'hC;
    Number6[16][14] = 4'hC;
    Number6[17][14] = 4'hF;
    Number6[18][14] = 4'hF;
    Number6[19][14] = 4'hF;
    Number6[20][14] = 4'hF;
    Number6[21][14] = 4'hF;
    Number6[22][14] = 4'hF;
    Number6[23][14] = 4'hF;
    Number6[0][15] = 4'hF;
    Number6[1][15] = 4'hF;
    Number6[2][15] = 4'hC;
    Number6[3][15] = 4'hC;
    Number6[4][15] = 4'hC;
    Number6[5][15] = 4'hC;
    Number6[6][15] = 4'hC;
    Number6[7][15] = 4'hC;
    Number6[8][15] = 4'hC;
    Number6[9][15] = 4'hC;
    Number6[10][15] = 4'hC;
    Number6[11][15] = 4'hC;
    Number6[12][15] = 4'hC;
    Number6[13][15] = 4'hC;
    Number6[14][15] = 4'hC;
    Number6[15][15] = 4'hC;
    Number6[16][15] = 4'hC;
    Number6[17][15] = 4'hF;
    Number6[18][15] = 4'hF;
    Number6[19][15] = 4'hF;
    Number6[20][15] = 4'hF;
    Number6[21][15] = 4'hF;
    Number6[22][15] = 4'hF;
    Number6[23][15] = 4'hF;
    Number6[0][16] = 4'hF;
    Number6[1][16] = 4'hF;
    Number6[2][16] = 4'hC;
    Number6[3][16] = 4'hC;
    Number6[4][16] = 4'hC;
    Number6[5][16] = 4'hC;
    Number6[6][16] = 4'hC;
    Number6[7][16] = 4'hC;
    Number6[8][16] = 4'hC;
    Number6[9][16] = 4'hC;
    Number6[10][16] = 4'hC;
    Number6[11][16] = 4'hC;
    Number6[12][16] = 4'hC;
    Number6[13][16] = 4'hC;
    Number6[14][16] = 4'hC;
    Number6[15][16] = 4'hC;
    Number6[16][16] = 4'hC;
    Number6[17][16] = 4'hF;
    Number6[18][16] = 4'hF;
    Number6[19][16] = 4'hF;
    Number6[20][16] = 4'hF;
    Number6[21][16] = 4'hF;
    Number6[22][16] = 4'hF;
    Number6[23][16] = 4'hF;
    Number6[0][17] = 4'hF;
    Number6[1][17] = 4'hF;
    Number6[2][17] = 4'hC;
    Number6[3][17] = 4'hC;
    Number6[4][17] = 4'hC;
    Number6[5][17] = 4'hC;
    Number6[6][17] = 4'hC;
    Number6[7][17] = 4'hC;
    Number6[8][17] = 4'hC;
    Number6[9][17] = 4'hC;
    Number6[10][17] = 4'hC;
    Number6[11][17] = 4'hC;
    Number6[12][17] = 4'hC;
    Number6[13][17] = 4'hC;
    Number6[14][17] = 4'hC;
    Number6[15][17] = 4'hC;
    Number6[16][17] = 4'hC;
    Number6[17][17] = 4'hF;
    Number6[18][17] = 4'hF;
    Number6[19][17] = 4'hF;
    Number6[20][17] = 4'hF;
    Number6[21][17] = 4'hF;
    Number6[22][17] = 4'hF;
    Number6[23][17] = 4'hF;
    Number6[0][18] = 4'hF;
    Number6[1][18] = 4'hF;
    Number6[2][18] = 4'hC;
    Number6[3][18] = 4'hC;
    Number6[4][18] = 4'hC;
    Number6[5][18] = 4'hC;
    Number6[6][18] = 4'hC;
    Number6[7][18] = 4'hF;
    Number6[8][18] = 4'hF;
    Number6[9][18] = 4'hF;
    Number6[10][18] = 4'hF;
    Number6[11][18] = 4'hF;
    Number6[12][18] = 4'hF;
    Number6[13][18] = 4'hF;
    Number6[14][18] = 4'hF;
    Number6[15][18] = 4'hF;
    Number6[16][18] = 4'hF;
    Number6[17][18] = 4'hC;
    Number6[18][18] = 4'hC;
    Number6[19][18] = 4'hC;
    Number6[20][18] = 4'hC;
    Number6[21][18] = 4'hC;
    Number6[22][18] = 4'hF;
    Number6[23][18] = 4'hF;
    Number6[0][19] = 4'hF;
    Number6[1][19] = 4'hF;
    Number6[2][19] = 4'hC;
    Number6[3][19] = 4'hC;
    Number6[4][19] = 4'hC;
    Number6[5][19] = 4'hC;
    Number6[6][19] = 4'hC;
    Number6[7][19] = 4'hF;
    Number6[8][19] = 4'hF;
    Number6[9][19] = 4'hF;
    Number6[10][19] = 4'hF;
    Number6[11][19] = 4'hF;
    Number6[12][19] = 4'hF;
    Number6[13][19] = 4'hF;
    Number6[14][19] = 4'hF;
    Number6[15][19] = 4'hF;
    Number6[16][19] = 4'hF;
    Number6[17][19] = 4'hC;
    Number6[18][19] = 4'hC;
    Number6[19][19] = 4'hC;
    Number6[20][19] = 4'hC;
    Number6[21][19] = 4'hC;
    Number6[22][19] = 4'hF;
    Number6[23][19] = 4'hF;
    Number6[0][20] = 4'hF;
    Number6[1][20] = 4'hF;
    Number6[2][20] = 4'hC;
    Number6[3][20] = 4'hC;
    Number6[4][20] = 4'hC;
    Number6[5][20] = 4'hC;
    Number6[6][20] = 4'hC;
    Number6[7][20] = 4'hF;
    Number6[8][20] = 4'hF;
    Number6[9][20] = 4'hF;
    Number6[10][20] = 4'hF;
    Number6[11][20] = 4'hF;
    Number6[12][20] = 4'hF;
    Number6[13][20] = 4'hF;
    Number6[14][20] = 4'hF;
    Number6[15][20] = 4'hF;
    Number6[16][20] = 4'hF;
    Number6[17][20] = 4'hC;
    Number6[18][20] = 4'hC;
    Number6[19][20] = 4'hC;
    Number6[20][20] = 4'hC;
    Number6[21][20] = 4'hC;
    Number6[22][20] = 4'hF;
    Number6[23][20] = 4'hF;
    Number6[0][21] = 4'hF;
    Number6[1][21] = 4'hF;
    Number6[2][21] = 4'hC;
    Number6[3][21] = 4'hC;
    Number6[4][21] = 4'hC;
    Number6[5][21] = 4'hC;
    Number6[6][21] = 4'hC;
    Number6[7][21] = 4'hF;
    Number6[8][21] = 4'hF;
    Number6[9][21] = 4'hF;
    Number6[10][21] = 4'hF;
    Number6[11][21] = 4'hF;
    Number6[12][21] = 4'hF;
    Number6[13][21] = 4'hF;
    Number6[14][21] = 4'hF;
    Number6[15][21] = 4'hF;
    Number6[16][21] = 4'hF;
    Number6[17][21] = 4'hC;
    Number6[18][21] = 4'hC;
    Number6[19][21] = 4'hC;
    Number6[20][21] = 4'hC;
    Number6[21][21] = 4'hC;
    Number6[22][21] = 4'hF;
    Number6[23][21] = 4'hF;
    Number6[0][22] = 4'hF;
    Number6[1][22] = 4'hF;
    Number6[2][22] = 4'hC;
    Number6[3][22] = 4'hC;
    Number6[4][22] = 4'hC;
    Number6[5][22] = 4'hC;
    Number6[6][22] = 4'hC;
    Number6[7][22] = 4'hF;
    Number6[8][22] = 4'hF;
    Number6[9][22] = 4'hF;
    Number6[10][22] = 4'hF;
    Number6[11][22] = 4'hF;
    Number6[12][22] = 4'hF;
    Number6[13][22] = 4'hF;
    Number6[14][22] = 4'hF;
    Number6[15][22] = 4'hF;
    Number6[16][22] = 4'hF;
    Number6[17][22] = 4'hC;
    Number6[18][22] = 4'hC;
    Number6[19][22] = 4'hC;
    Number6[20][22] = 4'hC;
    Number6[21][22] = 4'hC;
    Number6[22][22] = 4'hF;
    Number6[23][22] = 4'hF;
    Number6[0][23] = 4'hF;
    Number6[1][23] = 4'hF;
    Number6[2][23] = 4'hF;
    Number6[3][23] = 4'hF;
    Number6[4][23] = 4'hF;
    Number6[5][23] = 4'hF;
    Number6[6][23] = 4'hF;
    Number6[7][23] = 4'hC;
    Number6[8][23] = 4'hC;
    Number6[9][23] = 4'hC;
    Number6[10][23] = 4'hC;
    Number6[11][23] = 4'hC;
    Number6[12][23] = 4'hC;
    Number6[13][23] = 4'hC;
    Number6[14][23] = 4'hC;
    Number6[15][23] = 4'hC;
    Number6[16][23] = 4'hC;
    Number6[17][23] = 4'hF;
    Number6[18][23] = 4'hF;
    Number6[19][23] = 4'hF;
    Number6[20][23] = 4'hF;
    Number6[21][23] = 4'hF;
    Number6[22][23] = 4'hF;
    Number6[23][23] = 4'hF;
    Number6[0][24] = 4'hF;
    Number6[1][24] = 4'hF;
    Number6[2][24] = 4'hF;
    Number6[3][24] = 4'hF;
    Number6[4][24] = 4'hF;
    Number6[5][24] = 4'hF;
    Number6[6][24] = 4'hF;
    Number6[7][24] = 4'hC;
    Number6[8][24] = 4'hC;
    Number6[9][24] = 4'hC;
    Number6[10][24] = 4'hC;
    Number6[11][24] = 4'hC;
    Number6[12][24] = 4'hC;
    Number6[13][24] = 4'hC;
    Number6[14][24] = 4'hC;
    Number6[15][24] = 4'hC;
    Number6[16][24] = 4'hC;
    Number6[17][24] = 4'hF;
    Number6[18][24] = 4'hF;
    Number6[19][24] = 4'hF;
    Number6[20][24] = 4'hF;
    Number6[21][24] = 4'hF;
    Number6[22][24] = 4'hF;
    Number6[23][24] = 4'hF;
    Number6[0][25] = 4'hF;
    Number6[1][25] = 4'hF;
    Number6[2][25] = 4'hF;
    Number6[3][25] = 4'hF;
    Number6[4][25] = 4'hF;
    Number6[5][25] = 4'hF;
    Number6[6][25] = 4'hF;
    Number6[7][25] = 4'hC;
    Number6[8][25] = 4'hC;
    Number6[9][25] = 4'hC;
    Number6[10][25] = 4'hC;
    Number6[11][25] = 4'hC;
    Number6[12][25] = 4'hC;
    Number6[13][25] = 4'hC;
    Number6[14][25] = 4'hC;
    Number6[15][25] = 4'hC;
    Number6[16][25] = 4'hC;
    Number6[17][25] = 4'hF;
    Number6[18][25] = 4'hF;
    Number6[19][25] = 4'hF;
    Number6[20][25] = 4'hF;
    Number6[21][25] = 4'hF;
    Number6[22][25] = 4'hF;
    Number6[23][25] = 4'hF;
    Number6[0][26] = 4'hF;
    Number6[1][26] = 4'hF;
    Number6[2][26] = 4'hF;
    Number6[3][26] = 4'hF;
    Number6[4][26] = 4'hF;
    Number6[5][26] = 4'hF;
    Number6[6][26] = 4'hF;
    Number6[7][26] = 4'hC;
    Number6[8][26] = 4'hC;
    Number6[9][26] = 4'hC;
    Number6[10][26] = 4'hC;
    Number6[11][26] = 4'hC;
    Number6[12][26] = 4'hC;
    Number6[13][26] = 4'hC;
    Number6[14][26] = 4'hC;
    Number6[15][26] = 4'hC;
    Number6[16][26] = 4'hC;
    Number6[17][26] = 4'hF;
    Number6[18][26] = 4'hF;
    Number6[19][26] = 4'hF;
    Number6[20][26] = 4'hF;
    Number6[21][26] = 4'hF;
    Number6[22][26] = 4'hF;
    Number6[23][26] = 4'hF;
    Number6[0][27] = 4'hF;
    Number6[1][27] = 4'hF;
    Number6[2][27] = 4'hF;
    Number6[3][27] = 4'hF;
    Number6[4][27] = 4'hF;
    Number6[5][27] = 4'hF;
    Number6[6][27] = 4'hF;
    Number6[7][27] = 4'hC;
    Number6[8][27] = 4'hC;
    Number6[9][27] = 4'hC;
    Number6[10][27] = 4'hC;
    Number6[11][27] = 4'hC;
    Number6[12][27] = 4'hC;
    Number6[13][27] = 4'hC;
    Number6[14][27] = 4'hC;
    Number6[15][27] = 4'hC;
    Number6[16][27] = 4'hC;
    Number6[17][27] = 4'hF;
    Number6[18][27] = 4'hF;
    Number6[19][27] = 4'hF;
    Number6[20][27] = 4'hF;
    Number6[21][27] = 4'hF;
    Number6[22][27] = 4'hF;
    Number6[23][27] = 4'hF;
    Number6[0][28] = 4'hF;
    Number6[1][28] = 4'hF;
    Number6[2][28] = 4'hF;
    Number6[3][28] = 4'hF;
    Number6[4][28] = 4'hF;
    Number6[5][28] = 4'hF;
    Number6[6][28] = 4'hF;
    Number6[7][28] = 4'hF;
    Number6[8][28] = 4'hF;
    Number6[9][28] = 4'hF;
    Number6[10][28] = 4'hF;
    Number6[11][28] = 4'hF;
    Number6[12][28] = 4'hF;
    Number6[13][28] = 4'hF;
    Number6[14][28] = 4'hF;
    Number6[15][28] = 4'hF;
    Number6[16][28] = 4'hF;
    Number6[17][28] = 4'hF;
    Number6[18][28] = 4'hF;
    Number6[19][28] = 4'hF;
    Number6[20][28] = 4'hF;
    Number6[21][28] = 4'hF;
    Number6[22][28] = 4'hF;
    Number6[23][28] = 4'hF;
    Number6[0][29] = 4'hF;
    Number6[1][29] = 4'hF;
    Number6[2][29] = 4'hF;
    Number6[3][29] = 4'hF;
    Number6[4][29] = 4'hF;
    Number6[5][29] = 4'hF;
    Number6[6][29] = 4'hF;
    Number6[7][29] = 4'hF;
    Number6[8][29] = 4'hF;
    Number6[9][29] = 4'hF;
    Number6[10][29] = 4'hF;
    Number6[11][29] = 4'hF;
    Number6[12][29] = 4'hF;
    Number6[13][29] = 4'hF;
    Number6[14][29] = 4'hF;
    Number6[15][29] = 4'hF;
    Number6[16][29] = 4'hF;
    Number6[17][29] = 4'hF;
    Number6[18][29] = 4'hF;
    Number6[19][29] = 4'hF;
    Number6[20][29] = 4'hF;
    Number6[21][29] = 4'hF;
    Number6[22][29] = 4'hF;
    Number6[23][29] = 4'hF;
 
//Number 7
    Number7[0][0] = 4'hF;
    Number7[1][0] = 4'hF;
    Number7[2][0] = 4'hF;
    Number7[3][0] = 4'hF;
    Number7[4][0] = 4'hF;
    Number7[5][0] = 4'hF;
    Number7[6][0] = 4'hF;
    Number7[7][0] = 4'hF;
    Number7[8][0] = 4'hF;
    Number7[9][0] = 4'hF;
    Number7[10][0] = 4'hF;
    Number7[11][0] = 4'hF;
    Number7[12][0] = 4'hF;
    Number7[13][0] = 4'hF;
    Number7[14][0] = 4'hF;
    Number7[15][0] = 4'hF;
    Number7[16][0] = 4'hF;
    Number7[17][0] = 4'hF;
    Number7[18][0] = 4'hF;
    Number7[19][0] = 4'hF;
    Number7[20][0] = 4'hF;
    Number7[21][0] = 4'hF;
    Number7[22][0] = 4'hF;
    Number7[23][0] = 4'hF;
    Number7[0][1] = 4'hF;
    Number7[1][1] = 4'hF;
    Number7[2][1] = 4'hF;
    Number7[3][1] = 4'hF;
    Number7[4][1] = 4'hF;
    Number7[5][1] = 4'hF;
    Number7[6][1] = 4'hF;
    Number7[7][1] = 4'hF;
    Number7[8][1] = 4'hF;
    Number7[9][1] = 4'hF;
    Number7[10][1] = 4'hF;
    Number7[11][1] = 4'hF;
    Number7[12][1] = 4'hF;
    Number7[13][1] = 4'hF;
    Number7[14][1] = 4'hF;
    Number7[15][1] = 4'hF;
    Number7[16][1] = 4'hF;
    Number7[17][1] = 4'hF;
    Number7[18][1] = 4'hF;
    Number7[19][1] = 4'hF;
    Number7[20][1] = 4'hF;
    Number7[21][1] = 4'hF;
    Number7[22][1] = 4'hF;
    Number7[23][1] = 4'hF;
    Number7[0][2] = 4'hF;
    Number7[1][2] = 4'hF;
    Number7[2][2] = 4'hF;
    Number7[3][2] = 4'hF;
    Number7[4][2] = 4'hF;
    Number7[5][2] = 4'hF;
    Number7[6][2] = 4'hF;
    Number7[7][2] = 4'hF;
    Number7[8][2] = 4'hF;
    Number7[9][2] = 4'hF;
    Number7[10][2] = 4'hF;
    Number7[11][2] = 4'hF;
    Number7[12][2] = 4'hF;
    Number7[13][2] = 4'hF;
    Number7[14][2] = 4'hF;
    Number7[15][2] = 4'hF;
    Number7[16][2] = 4'hF;
    Number7[17][2] = 4'hF;
    Number7[18][2] = 4'hF;
    Number7[19][2] = 4'hF;
    Number7[20][2] = 4'hF;
    Number7[21][2] = 4'hF;
    Number7[22][2] = 4'hF;
    Number7[23][2] = 4'hF;
    Number7[0][3] = 4'hF;
    Number7[1][3] = 4'hF;
    Number7[2][3] = 4'hC;
    Number7[3][3] = 4'hC;
    Number7[4][3] = 4'hC;
    Number7[5][3] = 4'hC;
    Number7[6][3] = 4'hC;
    Number7[7][3] = 4'hC;
    Number7[8][3] = 4'hC;
    Number7[9][3] = 4'hC;
    Number7[10][3] = 4'hC;
    Number7[11][3] = 4'hC;
    Number7[12][3] = 4'hC;
    Number7[13][3] = 4'hC;
    Number7[14][3] = 4'hC;
    Number7[15][3] = 4'hC;
    Number7[16][3] = 4'hC;
    Number7[17][3] = 4'hC;
    Number7[18][3] = 4'hC;
    Number7[19][3] = 4'hC;
    Number7[20][3] = 4'hC;
    Number7[21][3] = 4'hC;
    Number7[22][3] = 4'hF;
    Number7[23][3] = 4'hF;
    Number7[0][4] = 4'hF;
    Number7[1][4] = 4'hF;
    Number7[2][4] = 4'hC;
    Number7[3][4] = 4'hC;
    Number7[4][4] = 4'hC;
    Number7[5][4] = 4'hC;
    Number7[6][4] = 4'hC;
    Number7[7][4] = 4'hC;
    Number7[8][4] = 4'hC;
    Number7[9][4] = 4'hC;
    Number7[10][4] = 4'hC;
    Number7[11][4] = 4'hC;
    Number7[12][4] = 4'hC;
    Number7[13][4] = 4'hC;
    Number7[14][4] = 4'hC;
    Number7[15][4] = 4'hC;
    Number7[16][4] = 4'hC;
    Number7[17][4] = 4'hC;
    Number7[18][4] = 4'hC;
    Number7[19][4] = 4'hC;
    Number7[20][4] = 4'hC;
    Number7[21][4] = 4'hC;
    Number7[22][4] = 4'hF;
    Number7[23][4] = 4'hF;
    Number7[0][5] = 4'hF;
    Number7[1][5] = 4'hF;
    Number7[2][5] = 4'hC;
    Number7[3][5] = 4'hC;
    Number7[4][5] = 4'hC;
    Number7[5][5] = 4'hC;
    Number7[6][5] = 4'hC;
    Number7[7][5] = 4'hC;
    Number7[8][5] = 4'hC;
    Number7[9][5] = 4'hC;
    Number7[10][5] = 4'hC;
    Number7[11][5] = 4'hC;
    Number7[12][5] = 4'hC;
    Number7[13][5] = 4'hC;
    Number7[14][5] = 4'hC;
    Number7[15][5] = 4'hC;
    Number7[16][5] = 4'hC;
    Number7[17][5] = 4'hC;
    Number7[18][5] = 4'hC;
    Number7[19][5] = 4'hC;
    Number7[20][5] = 4'hC;
    Number7[21][5] = 4'hC;
    Number7[22][5] = 4'hF;
    Number7[23][5] = 4'hF;
    Number7[0][6] = 4'hF;
    Number7[1][6] = 4'hF;
    Number7[2][6] = 4'hC;
    Number7[3][6] = 4'hC;
    Number7[4][6] = 4'hC;
    Number7[5][6] = 4'hC;
    Number7[6][6] = 4'hC;
    Number7[7][6] = 4'hC;
    Number7[8][6] = 4'hC;
    Number7[9][6] = 4'hC;
    Number7[10][6] = 4'hC;
    Number7[11][6] = 4'hC;
    Number7[12][6] = 4'hC;
    Number7[13][6] = 4'hC;
    Number7[14][6] = 4'hC;
    Number7[15][6] = 4'hC;
    Number7[16][6] = 4'hC;
    Number7[17][6] = 4'hC;
    Number7[18][6] = 4'hC;
    Number7[19][6] = 4'hC;
    Number7[20][6] = 4'hC;
    Number7[21][6] = 4'hC;
    Number7[22][6] = 4'hF;
    Number7[23][6] = 4'hF;
    Number7[0][7] = 4'hF;
    Number7[1][7] = 4'hF;
    Number7[2][7] = 4'hC;
    Number7[3][7] = 4'hC;
    Number7[4][7] = 4'hC;
    Number7[5][7] = 4'hC;
    Number7[6][7] = 4'hC;
    Number7[7][7] = 4'hC;
    Number7[8][7] = 4'hC;
    Number7[9][7] = 4'hC;
    Number7[10][7] = 4'hC;
    Number7[11][7] = 4'hC;
    Number7[12][7] = 4'hC;
    Number7[13][7] = 4'hC;
    Number7[14][7] = 4'hC;
    Number7[15][7] = 4'hC;
    Number7[16][7] = 4'hC;
    Number7[17][7] = 4'hC;
    Number7[18][7] = 4'hC;
    Number7[19][7] = 4'hC;
    Number7[20][7] = 4'hC;
    Number7[21][7] = 4'hC;
    Number7[22][7] = 4'hF;
    Number7[23][7] = 4'hF;
    Number7[0][8] = 4'hF;
    Number7[1][8] = 4'hF;
    Number7[2][8] = 4'hF;
    Number7[3][8] = 4'hF;
    Number7[4][8] = 4'hF;
    Number7[5][8] = 4'hF;
    Number7[6][8] = 4'hF;
    Number7[7][8] = 4'hF;
    Number7[8][8] = 4'hF;
    Number7[9][8] = 4'hF;
    Number7[10][8] = 4'hF;
    Number7[11][8] = 4'hF;
    Number7[12][8] = 4'hF;
    Number7[13][8] = 4'hF;
    Number7[14][8] = 4'hF;
    Number7[15][8] = 4'hF;
    Number7[16][8] = 4'hF;
    Number7[17][8] = 4'hC;
    Number7[18][8] = 4'hC;
    Number7[19][8] = 4'hC;
    Number7[20][8] = 4'hC;
    Number7[21][8] = 4'hC;
    Number7[22][8] = 4'hF;
    Number7[23][8] = 4'hF;
    Number7[0][9] = 4'hF;
    Number7[1][9] = 4'hF;
    Number7[2][9] = 4'hF;
    Number7[3][9] = 4'hF;
    Number7[4][9] = 4'hF;
    Number7[5][9] = 4'hF;
    Number7[6][9] = 4'hF;
    Number7[7][9] = 4'hF;
    Number7[8][9] = 4'hF;
    Number7[9][9] = 4'hF;
    Number7[10][9] = 4'hF;
    Number7[11][9] = 4'hF;
    Number7[12][9] = 4'hF;
    Number7[13][9] = 4'hF;
    Number7[14][9] = 4'hF;
    Number7[15][9] = 4'hF;
    Number7[16][9] = 4'hF;
    Number7[17][9] = 4'hC;
    Number7[18][9] = 4'hC;
    Number7[19][9] = 4'hC;
    Number7[20][9] = 4'hC;
    Number7[21][9] = 4'hC;
    Number7[22][9] = 4'hF;
    Number7[23][9] = 4'hF;
    Number7[0][10] = 4'hF;
    Number7[1][10] = 4'hF;
    Number7[2][10] = 4'hF;
    Number7[3][10] = 4'hF;
    Number7[4][10] = 4'hF;
    Number7[5][10] = 4'hF;
    Number7[6][10] = 4'hF;
    Number7[7][10] = 4'hF;
    Number7[8][10] = 4'hF;
    Number7[9][10] = 4'hF;
    Number7[10][10] = 4'hF;
    Number7[11][10] = 4'hF;
    Number7[12][10] = 4'hF;
    Number7[13][10] = 4'hF;
    Number7[14][10] = 4'hF;
    Number7[15][10] = 4'hF;
    Number7[16][10] = 4'hF;
    Number7[17][10] = 4'hC;
    Number7[18][10] = 4'hC;
    Number7[19][10] = 4'hC;
    Number7[20][10] = 4'hC;
    Number7[21][10] = 4'hC;
    Number7[22][10] = 4'hF;
    Number7[23][10] = 4'hF;
    Number7[0][11] = 4'hF;
    Number7[1][11] = 4'hF;
    Number7[2][11] = 4'hF;
    Number7[3][11] = 4'hF;
    Number7[4][11] = 4'hF;
    Number7[5][11] = 4'hF;
    Number7[6][11] = 4'hF;
    Number7[7][11] = 4'hF;
    Number7[8][11] = 4'hF;
    Number7[9][11] = 4'hF;
    Number7[10][11] = 4'hF;
    Number7[11][11] = 4'hF;
    Number7[12][11] = 4'hF;
    Number7[13][11] = 4'hF;
    Number7[14][11] = 4'hF;
    Number7[15][11] = 4'hF;
    Number7[16][11] = 4'hF;
    Number7[17][11] = 4'hC;
    Number7[18][11] = 4'hC;
    Number7[19][11] = 4'hC;
    Number7[20][11] = 4'hC;
    Number7[21][11] = 4'hC;
    Number7[22][11] = 4'hF;
    Number7[23][11] = 4'hF;
    Number7[0][12] = 4'hF;
    Number7[1][12] = 4'hF;
    Number7[2][12] = 4'hF;
    Number7[3][12] = 4'hF;
    Number7[4][12] = 4'hF;
    Number7[5][12] = 4'hF;
    Number7[6][12] = 4'hF;
    Number7[7][12] = 4'hF;
    Number7[8][12] = 4'hF;
    Number7[9][12] = 4'hF;
    Number7[10][12] = 4'hF;
    Number7[11][12] = 4'hF;
    Number7[12][12] = 4'hF;
    Number7[13][12] = 4'hF;
    Number7[14][12] = 4'hF;
    Number7[15][12] = 4'hF;
    Number7[16][12] = 4'hF;
    Number7[17][12] = 4'hC;
    Number7[18][12] = 4'hC;
    Number7[19][12] = 4'hC;
    Number7[20][12] = 4'hC;
    Number7[21][12] = 4'hC;
    Number7[22][12] = 4'hF;
    Number7[23][12] = 4'hF;
    Number7[0][13] = 4'hF;
    Number7[1][13] = 4'hF;
    Number7[2][13] = 4'hF;
    Number7[3][13] = 4'hF;
    Number7[4][13] = 4'hF;
    Number7[5][13] = 4'hF;
    Number7[6][13] = 4'hF;
    Number7[7][13] = 4'hF;
    Number7[8][13] = 4'hF;
    Number7[9][13] = 4'hF;
    Number7[10][13] = 4'hF;
    Number7[11][13] = 4'hF;
    Number7[12][13] = 4'hC;
    Number7[13][13] = 4'hC;
    Number7[14][13] = 4'hC;
    Number7[15][13] = 4'hC;
    Number7[16][13] = 4'hC;
    Number7[17][13] = 4'hF;
    Number7[18][13] = 4'hF;
    Number7[19][13] = 4'hF;
    Number7[20][13] = 4'hF;
    Number7[21][13] = 4'hF;
    Number7[22][13] = 4'hF;
    Number7[23][13] = 4'hF;
    Number7[0][14] = 4'hF;
    Number7[1][14] = 4'hF;
    Number7[2][14] = 4'hF;
    Number7[3][14] = 4'hF;
    Number7[4][14] = 4'hF;
    Number7[5][14] = 4'hF;
    Number7[6][14] = 4'hF;
    Number7[7][14] = 4'hF;
    Number7[8][14] = 4'hF;
    Number7[9][14] = 4'hF;
    Number7[10][14] = 4'hF;
    Number7[11][14] = 4'hF;
    Number7[12][14] = 4'hC;
    Number7[13][14] = 4'hC;
    Number7[14][14] = 4'hC;
    Number7[15][14] = 4'hC;
    Number7[16][14] = 4'hC;
    Number7[17][14] = 4'hF;
    Number7[18][14] = 4'hF;
    Number7[19][14] = 4'hF;
    Number7[20][14] = 4'hF;
    Number7[21][14] = 4'hF;
    Number7[22][14] = 4'hF;
    Number7[23][14] = 4'hF;
    Number7[0][15] = 4'hF;
    Number7[1][15] = 4'hF;
    Number7[2][15] = 4'hF;
    Number7[3][15] = 4'hF;
    Number7[4][15] = 4'hF;
    Number7[5][15] = 4'hF;
    Number7[6][15] = 4'hF;
    Number7[7][15] = 4'hF;
    Number7[8][15] = 4'hF;
    Number7[9][15] = 4'hF;
    Number7[10][15] = 4'hF;
    Number7[11][15] = 4'hF;
    Number7[12][15] = 4'hC;
    Number7[13][15] = 4'hC;
    Number7[14][15] = 4'hC;
    Number7[15][15] = 4'hC;
    Number7[16][15] = 4'hC;
    Number7[17][15] = 4'hF;
    Number7[18][15] = 4'hF;
    Number7[19][15] = 4'hF;
    Number7[20][15] = 4'hF;
    Number7[21][15] = 4'hF;
    Number7[22][15] = 4'hF;
    Number7[23][15] = 4'hF;
    Number7[0][16] = 4'hF;
    Number7[1][16] = 4'hF;
    Number7[2][16] = 4'hF;
    Number7[3][16] = 4'hF;
    Number7[4][16] = 4'hF;
    Number7[5][16] = 4'hF;
    Number7[6][16] = 4'hF;
    Number7[7][16] = 4'hF;
    Number7[8][16] = 4'hF;
    Number7[9][16] = 4'hF;
    Number7[10][16] = 4'hF;
    Number7[11][16] = 4'hF;
    Number7[12][16] = 4'hC;
    Number7[13][16] = 4'hC;
    Number7[14][16] = 4'hC;
    Number7[15][16] = 4'hC;
    Number7[16][16] = 4'hC;
    Number7[17][16] = 4'hF;
    Number7[18][16] = 4'hF;
    Number7[19][16] = 4'hF;
    Number7[20][16] = 4'hF;
    Number7[21][16] = 4'hF;
    Number7[22][16] = 4'hF;
    Number7[23][16] = 4'hF;
    Number7[0][17] = 4'hF;
    Number7[1][17] = 4'hF;
    Number7[2][17] = 4'hF;
    Number7[3][17] = 4'hF;
    Number7[4][17] = 4'hF;
    Number7[5][17] = 4'hF;
    Number7[6][17] = 4'hF;
    Number7[7][17] = 4'hF;
    Number7[8][17] = 4'hF;
    Number7[9][17] = 4'hF;
    Number7[10][17] = 4'hF;
    Number7[11][17] = 4'hF;
    Number7[12][17] = 4'hC;
    Number7[13][17] = 4'hC;
    Number7[14][17] = 4'hC;
    Number7[15][17] = 4'hC;
    Number7[16][17] = 4'hC;
    Number7[17][17] = 4'hF;
    Number7[18][17] = 4'hF;
    Number7[19][17] = 4'hF;
    Number7[20][17] = 4'hF;
    Number7[21][17] = 4'hF;
    Number7[22][17] = 4'hF;
    Number7[23][17] = 4'hF;
    Number7[0][18] = 4'hF;
    Number7[1][18] = 4'hF;
    Number7[2][18] = 4'hF;
    Number7[3][18] = 4'hF;
    Number7[4][18] = 4'hF;
    Number7[5][18] = 4'hF;
    Number7[6][18] = 4'hF;
    Number7[7][18] = 4'hC;
    Number7[8][18] = 4'hC;
    Number7[9][18] = 4'hC;
    Number7[10][18] = 4'hC;
    Number7[11][18] = 4'hC;
    Number7[12][18] = 4'hF;
    Number7[13][18] = 4'hF;
    Number7[14][18] = 4'hF;
    Number7[15][18] = 4'hF;
    Number7[16][18] = 4'hF;
    Number7[17][18] = 4'hF;
    Number7[18][18] = 4'hF;
    Number7[19][18] = 4'hF;
    Number7[20][18] = 4'hF;
    Number7[21][18] = 4'hF;
    Number7[22][18] = 4'hF;
    Number7[23][18] = 4'hF;
    Number7[0][19] = 4'hF;
    Number7[1][19] = 4'hF;
    Number7[2][19] = 4'hF;
    Number7[3][19] = 4'hF;
    Number7[4][19] = 4'hF;
    Number7[5][19] = 4'hF;
    Number7[6][19] = 4'hF;
    Number7[7][19] = 4'hC;
    Number7[8][19] = 4'hC;
    Number7[9][19] = 4'hC;
    Number7[10][19] = 4'hC;
    Number7[11][19] = 4'hC;
    Number7[12][19] = 4'hF;
    Number7[13][19] = 4'hF;
    Number7[14][19] = 4'hF;
    Number7[15][19] = 4'hF;
    Number7[16][19] = 4'hF;
    Number7[17][19] = 4'hF;
    Number7[18][19] = 4'hF;
    Number7[19][19] = 4'hF;
    Number7[20][19] = 4'hF;
    Number7[21][19] = 4'hF;
    Number7[22][19] = 4'hF;
    Number7[23][19] = 4'hF;
    Number7[0][20] = 4'hF;
    Number7[1][20] = 4'hF;
    Number7[2][20] = 4'hF;
    Number7[3][20] = 4'hF;
    Number7[4][20] = 4'hF;
    Number7[5][20] = 4'hF;
    Number7[6][20] = 4'hF;
    Number7[7][20] = 4'hC;
    Number7[8][20] = 4'hC;
    Number7[9][20] = 4'hC;
    Number7[10][20] = 4'hC;
    Number7[11][20] = 4'hC;
    Number7[12][20] = 4'hF;
    Number7[13][20] = 4'hF;
    Number7[14][20] = 4'hF;
    Number7[15][20] = 4'hF;
    Number7[16][20] = 4'hF;
    Number7[17][20] = 4'hF;
    Number7[18][20] = 4'hF;
    Number7[19][20] = 4'hF;
    Number7[20][20] = 4'hF;
    Number7[21][20] = 4'hF;
    Number7[22][20] = 4'hF;
    Number7[23][20] = 4'hF;
    Number7[0][21] = 4'hF;
    Number7[1][21] = 4'hF;
    Number7[2][21] = 4'hF;
    Number7[3][21] = 4'hF;
    Number7[4][21] = 4'hF;
    Number7[5][21] = 4'hF;
    Number7[6][21] = 4'hF;
    Number7[7][21] = 4'hC;
    Number7[8][21] = 4'hC;
    Number7[9][21] = 4'hC;
    Number7[10][21] = 4'hC;
    Number7[11][21] = 4'hC;
    Number7[12][21] = 4'hF;
    Number7[13][21] = 4'hF;
    Number7[14][21] = 4'hF;
    Number7[15][21] = 4'hF;
    Number7[16][21] = 4'hF;
    Number7[17][21] = 4'hF;
    Number7[18][21] = 4'hF;
    Number7[19][21] = 4'hF;
    Number7[20][21] = 4'hF;
    Number7[21][21] = 4'hF;
    Number7[22][21] = 4'hF;
    Number7[23][21] = 4'hF;
    Number7[0][22] = 4'hF;
    Number7[1][22] = 4'hF;
    Number7[2][22] = 4'hF;
    Number7[3][22] = 4'hF;
    Number7[4][22] = 4'hF;
    Number7[5][22] = 4'hF;
    Number7[6][22] = 4'hF;
    Number7[7][22] = 4'hC;
    Number7[8][22] = 4'hC;
    Number7[9][22] = 4'hC;
    Number7[10][22] = 4'hC;
    Number7[11][22] = 4'hC;
    Number7[12][22] = 4'hF;
    Number7[13][22] = 4'hF;
    Number7[14][22] = 4'hF;
    Number7[15][22] = 4'hF;
    Number7[16][22] = 4'hF;
    Number7[17][22] = 4'hF;
    Number7[18][22] = 4'hF;
    Number7[19][22] = 4'hF;
    Number7[20][22] = 4'hF;
    Number7[21][22] = 4'hF;
    Number7[22][22] = 4'hF;
    Number7[23][22] = 4'hF;
    Number7[0][23] = 4'hF;
    Number7[1][23] = 4'hF;
    Number7[2][23] = 4'hF;
    Number7[3][23] = 4'hF;
    Number7[4][23] = 4'hF;
    Number7[5][23] = 4'hF;
    Number7[6][23] = 4'hF;
    Number7[7][23] = 4'hC;
    Number7[8][23] = 4'hC;
    Number7[9][23] = 4'hC;
    Number7[10][23] = 4'hC;
    Number7[11][23] = 4'hC;
    Number7[12][23] = 4'hF;
    Number7[13][23] = 4'hF;
    Number7[14][23] = 4'hF;
    Number7[15][23] = 4'hF;
    Number7[16][23] = 4'hF;
    Number7[17][23] = 4'hF;
    Number7[18][23] = 4'hF;
    Number7[19][23] = 4'hF;
    Number7[20][23] = 4'hF;
    Number7[21][23] = 4'hF;
    Number7[22][23] = 4'hF;
    Number7[23][23] = 4'hF;
    Number7[0][24] = 4'hF;
    Number7[1][24] = 4'hF;
    Number7[2][24] = 4'hF;
    Number7[3][24] = 4'hF;
    Number7[4][24] = 4'hF;
    Number7[5][24] = 4'hF;
    Number7[6][24] = 4'hF;
    Number7[7][24] = 4'hC;
    Number7[8][24] = 4'hC;
    Number7[9][24] = 4'hC;
    Number7[10][24] = 4'hC;
    Number7[11][24] = 4'hC;
    Number7[12][24] = 4'hF;
    Number7[13][24] = 4'hF;
    Number7[14][24] = 4'hF;
    Number7[15][24] = 4'hF;
    Number7[16][24] = 4'hF;
    Number7[17][24] = 4'hF;
    Number7[18][24] = 4'hF;
    Number7[19][24] = 4'hF;
    Number7[20][24] = 4'hF;
    Number7[21][24] = 4'hF;
    Number7[22][24] = 4'hF;
    Number7[23][24] = 4'hF;
    Number7[0][25] = 4'hF;
    Number7[1][25] = 4'hF;
    Number7[2][25] = 4'hF;
    Number7[3][25] = 4'hF;
    Number7[4][25] = 4'hF;
    Number7[5][25] = 4'hF;
    Number7[6][25] = 4'hF;
    Number7[7][25] = 4'hC;
    Number7[8][25] = 4'hC;
    Number7[9][25] = 4'hC;
    Number7[10][25] = 4'hC;
    Number7[11][25] = 4'hC;
    Number7[12][25] = 4'hF;
    Number7[13][25] = 4'hF;
    Number7[14][25] = 4'hF;
    Number7[15][25] = 4'hF;
    Number7[16][25] = 4'hF;
    Number7[17][25] = 4'hF;
    Number7[18][25] = 4'hF;
    Number7[19][25] = 4'hF;
    Number7[20][25] = 4'hF;
    Number7[21][25] = 4'hF;
    Number7[22][25] = 4'hF;
    Number7[23][25] = 4'hF;
    Number7[0][26] = 4'hF;
    Number7[1][26] = 4'hF;
    Number7[2][26] = 4'hF;
    Number7[3][26] = 4'hF;
    Number7[4][26] = 4'hF;
    Number7[5][26] = 4'hF;
    Number7[6][26] = 4'hF;
    Number7[7][26] = 4'hC;
    Number7[8][26] = 4'hC;
    Number7[9][26] = 4'hC;
    Number7[10][26] = 4'hC;
    Number7[11][26] = 4'hC;
    Number7[12][26] = 4'hF;
    Number7[13][26] = 4'hF;
    Number7[14][26] = 4'hF;
    Number7[15][26] = 4'hF;
    Number7[16][26] = 4'hF;
    Number7[17][26] = 4'hF;
    Number7[18][26] = 4'hF;
    Number7[19][26] = 4'hF;
    Number7[20][26] = 4'hF;
    Number7[21][26] = 4'hF;
    Number7[22][26] = 4'hF;
    Number7[23][26] = 4'hF;
    Number7[0][27] = 4'hF;
    Number7[1][27] = 4'hF;
    Number7[2][27] = 4'hF;
    Number7[3][27] = 4'hF;
    Number7[4][27] = 4'hF;
    Number7[5][27] = 4'hF;
    Number7[6][27] = 4'hF;
    Number7[7][27] = 4'hC;
    Number7[8][27] = 4'hC;
    Number7[9][27] = 4'hC;
    Number7[10][27] = 4'hC;
    Number7[11][27] = 4'hC;
    Number7[12][27] = 4'hF;
    Number7[13][27] = 4'hF;
    Number7[14][27] = 4'hF;
    Number7[15][27] = 4'hF;
    Number7[16][27] = 4'hF;
    Number7[17][27] = 4'hF;
    Number7[18][27] = 4'hF;
    Number7[19][27] = 4'hF;
    Number7[20][27] = 4'hF;
    Number7[21][27] = 4'hF;
    Number7[22][27] = 4'hF;
    Number7[23][27] = 4'hF;
    Number7[0][28] = 4'hF;
    Number7[1][28] = 4'hF;
    Number7[2][28] = 4'hF;
    Number7[3][28] = 4'hF;
    Number7[4][28] = 4'hF;
    Number7[5][28] = 4'hF;
    Number7[6][28] = 4'hF;
    Number7[7][28] = 4'hF;
    Number7[8][28] = 4'hF;
    Number7[9][28] = 4'hF;
    Number7[10][28] = 4'hF;
    Number7[11][28] = 4'hF;
    Number7[12][28] = 4'hF;
    Number7[13][28] = 4'hF;
    Number7[14][28] = 4'hF;
    Number7[15][28] = 4'hF;
    Number7[16][28] = 4'hF;
    Number7[17][28] = 4'hF;
    Number7[18][28] = 4'hF;
    Number7[19][28] = 4'hF;
    Number7[20][28] = 4'hF;
    Number7[21][28] = 4'hF;
    Number7[22][28] = 4'hF;
    Number7[23][28] = 4'hF;
    Number7[0][29] = 4'hF;
    Number7[1][29] = 4'hF;
    Number7[2][29] = 4'hF;
    Number7[3][29] = 4'hF;
    Number7[4][29] = 4'hF;
    Number7[5][29] = 4'hF;
    Number7[6][29] = 4'hF;
    Number7[7][29] = 4'hF;
    Number7[8][29] = 4'hF;
    Number7[9][29] = 4'hF;
    Number7[10][29] = 4'hF;
    Number7[11][29] = 4'hF;
    Number7[12][29] = 4'hF;
    Number7[13][29] = 4'hF;
    Number7[14][29] = 4'hF;
    Number7[15][29] = 4'hF;
    Number7[16][29] = 4'hF;
    Number7[17][29] = 4'hF;
    Number7[18][29] = 4'hF;
    Number7[19][29] = 4'hF;
    Number7[20][29] = 4'hF;
    Number7[21][29] = 4'hF;
    Number7[22][29] = 4'hF;
    Number7[23][29] = 4'hF;
 
//Number 8
    Number8[0][0] = 4'hF;
    Number8[1][0] = 4'hF;
    Number8[2][0] = 4'hF;
    Number8[3][0] = 4'hF;
    Number8[4][0] = 4'hF;
    Number8[5][0] = 4'hF;
    Number8[6][0] = 4'hF;
    Number8[7][0] = 4'hF;
    Number8[8][0] = 4'hF;
    Number8[9][0] = 4'hF;
    Number8[10][0] = 4'hF;
    Number8[11][0] = 4'hF;
    Number8[12][0] = 4'hF;
    Number8[13][0] = 4'hF;
    Number8[14][0] = 4'hF;
    Number8[15][0] = 4'hF;
    Number8[16][0] = 4'hF;
    Number8[17][0] = 4'hF;
    Number8[18][0] = 4'hF;
    Number8[19][0] = 4'hF;
    Number8[20][0] = 4'hF;
    Number8[21][0] = 4'hF;
    Number8[22][0] = 4'hF;
    Number8[23][0] = 4'hF;
    Number8[0][1] = 4'hF;
    Number8[1][1] = 4'hF;
    Number8[2][1] = 4'hF;
    Number8[3][1] = 4'hF;
    Number8[4][1] = 4'hF;
    Number8[5][1] = 4'hF;
    Number8[6][1] = 4'hF;
    Number8[7][1] = 4'hF;
    Number8[8][1] = 4'hF;
    Number8[9][1] = 4'hF;
    Number8[10][1] = 4'hF;
    Number8[11][1] = 4'hF;
    Number8[12][1] = 4'hF;
    Number8[13][1] = 4'hF;
    Number8[14][1] = 4'hF;
    Number8[15][1] = 4'hF;
    Number8[16][1] = 4'hF;
    Number8[17][1] = 4'hF;
    Number8[18][1] = 4'hF;
    Number8[19][1] = 4'hF;
    Number8[20][1] = 4'hF;
    Number8[21][1] = 4'hF;
    Number8[22][1] = 4'hF;
    Number8[23][1] = 4'hF;
    Number8[0][2] = 4'hF;
    Number8[1][2] = 4'hF;
    Number8[2][2] = 4'hF;
    Number8[3][2] = 4'hF;
    Number8[4][2] = 4'hF;
    Number8[5][2] = 4'hF;
    Number8[6][2] = 4'hF;
    Number8[7][2] = 4'hF;
    Number8[8][2] = 4'hF;
    Number8[9][2] = 4'hF;
    Number8[10][2] = 4'hF;
    Number8[11][2] = 4'hF;
    Number8[12][2] = 4'hF;
    Number8[13][2] = 4'hF;
    Number8[14][2] = 4'hF;
    Number8[15][2] = 4'hF;
    Number8[16][2] = 4'hF;
    Number8[17][2] = 4'hF;
    Number8[18][2] = 4'hF;
    Number8[19][2] = 4'hF;
    Number8[20][2] = 4'hF;
    Number8[21][2] = 4'hF;
    Number8[22][2] = 4'hF;
    Number8[23][2] = 4'hF;
    Number8[0][3] = 4'hF;
    Number8[1][3] = 4'hF;
    Number8[2][3] = 4'hF;
    Number8[3][3] = 4'hF;
    Number8[4][3] = 4'hF;
    Number8[5][3] = 4'hF;
    Number8[6][3] = 4'hF;
    Number8[7][3] = 4'hC;
    Number8[8][3] = 4'hC;
    Number8[9][3] = 4'hC;
    Number8[10][3] = 4'hC;
    Number8[11][3] = 4'hC;
    Number8[12][3] = 4'hC;
    Number8[13][3] = 4'hC;
    Number8[14][3] = 4'hC;
    Number8[15][3] = 4'hC;
    Number8[16][3] = 4'hC;
    Number8[17][3] = 4'hF;
    Number8[18][3] = 4'hF;
    Number8[19][3] = 4'hF;
    Number8[20][3] = 4'hF;
    Number8[21][3] = 4'hF;
    Number8[22][3] = 4'hF;
    Number8[23][3] = 4'hF;
    Number8[0][4] = 4'hF;
    Number8[1][4] = 4'hF;
    Number8[2][4] = 4'hF;
    Number8[3][4] = 4'hF;
    Number8[4][4] = 4'hF;
    Number8[5][4] = 4'hF;
    Number8[6][4] = 4'hF;
    Number8[7][4] = 4'hC;
    Number8[8][4] = 4'hC;
    Number8[9][4] = 4'hC;
    Number8[10][4] = 4'hC;
    Number8[11][4] = 4'hC;
    Number8[12][4] = 4'hC;
    Number8[13][4] = 4'hC;
    Number8[14][4] = 4'hC;
    Number8[15][4] = 4'hC;
    Number8[16][4] = 4'hC;
    Number8[17][4] = 4'hF;
    Number8[18][4] = 4'hF;
    Number8[19][4] = 4'hF;
    Number8[20][4] = 4'hF;
    Number8[21][4] = 4'hF;
    Number8[22][4] = 4'hF;
    Number8[23][4] = 4'hF;
    Number8[0][5] = 4'hF;
    Number8[1][5] = 4'hF;
    Number8[2][5] = 4'hF;
    Number8[3][5] = 4'hF;
    Number8[4][5] = 4'hF;
    Number8[5][5] = 4'hF;
    Number8[6][5] = 4'hF;
    Number8[7][5] = 4'hC;
    Number8[8][5] = 4'hC;
    Number8[9][5] = 4'hC;
    Number8[10][5] = 4'hC;
    Number8[11][5] = 4'hC;
    Number8[12][5] = 4'hC;
    Number8[13][5] = 4'hC;
    Number8[14][5] = 4'hC;
    Number8[15][5] = 4'hC;
    Number8[16][5] = 4'hC;
    Number8[17][5] = 4'hF;
    Number8[18][5] = 4'hF;
    Number8[19][5] = 4'hF;
    Number8[20][5] = 4'hF;
    Number8[21][5] = 4'hF;
    Number8[22][5] = 4'hF;
    Number8[23][5] = 4'hF;
    Number8[0][6] = 4'hF;
    Number8[1][6] = 4'hF;
    Number8[2][6] = 4'hF;
    Number8[3][6] = 4'hF;
    Number8[4][6] = 4'hF;
    Number8[5][6] = 4'hF;
    Number8[6][6] = 4'hF;
    Number8[7][6] = 4'hC;
    Number8[8][6] = 4'hC;
    Number8[9][6] = 4'hC;
    Number8[10][6] = 4'hC;
    Number8[11][6] = 4'hC;
    Number8[12][6] = 4'hC;
    Number8[13][6] = 4'hC;
    Number8[14][6] = 4'hC;
    Number8[15][6] = 4'hC;
    Number8[16][6] = 4'hC;
    Number8[17][6] = 4'hF;
    Number8[18][6] = 4'hF;
    Number8[19][6] = 4'hF;
    Number8[20][6] = 4'hF;
    Number8[21][6] = 4'hF;
    Number8[22][6] = 4'hF;
    Number8[23][6] = 4'hF;
    Number8[0][7] = 4'hF;
    Number8[1][7] = 4'hF;
    Number8[2][7] = 4'hF;
    Number8[3][7] = 4'hF;
    Number8[4][7] = 4'hF;
    Number8[5][7] = 4'hF;
    Number8[6][7] = 4'hF;
    Number8[7][7] = 4'hC;
    Number8[8][7] = 4'hC;
    Number8[9][7] = 4'hC;
    Number8[10][7] = 4'hC;
    Number8[11][7] = 4'hC;
    Number8[12][7] = 4'hC;
    Number8[13][7] = 4'hC;
    Number8[14][7] = 4'hC;
    Number8[15][7] = 4'hC;
    Number8[16][7] = 4'hC;
    Number8[17][7] = 4'hF;
    Number8[18][7] = 4'hF;
    Number8[19][7] = 4'hF;
    Number8[20][7] = 4'hF;
    Number8[21][7] = 4'hF;
    Number8[22][7] = 4'hF;
    Number8[23][7] = 4'hF;
    Number8[0][8] = 4'hF;
    Number8[1][8] = 4'hF;
    Number8[2][8] = 4'hC;
    Number8[3][8] = 4'hC;
    Number8[4][8] = 4'hC;
    Number8[5][8] = 4'hC;
    Number8[6][8] = 4'hC;
    Number8[7][8] = 4'hF;
    Number8[8][8] = 4'hF;
    Number8[9][8] = 4'hF;
    Number8[10][8] = 4'hF;
    Number8[11][8] = 4'hF;
    Number8[12][8] = 4'hF;
    Number8[13][8] = 4'hF;
    Number8[14][8] = 4'hF;
    Number8[15][8] = 4'hF;
    Number8[16][8] = 4'hF;
    Number8[17][8] = 4'hC;
    Number8[18][8] = 4'hC;
    Number8[19][8] = 4'hC;
    Number8[20][8] = 4'hC;
    Number8[21][8] = 4'hC;
    Number8[22][8] = 4'hF;
    Number8[23][8] = 4'hF;
    Number8[0][9] = 4'hF;
    Number8[1][9] = 4'hF;
    Number8[2][9] = 4'hC;
    Number8[3][9] = 4'hC;
    Number8[4][9] = 4'hC;
    Number8[5][9] = 4'hC;
    Number8[6][9] = 4'hC;
    Number8[7][9] = 4'hF;
    Number8[8][9] = 4'hF;
    Number8[9][9] = 4'hF;
    Number8[10][9] = 4'hF;
    Number8[11][9] = 4'hF;
    Number8[12][9] = 4'hF;
    Number8[13][9] = 4'hF;
    Number8[14][9] = 4'hF;
    Number8[15][9] = 4'hF;
    Number8[16][9] = 4'hF;
    Number8[17][9] = 4'hC;
    Number8[18][9] = 4'hC;
    Number8[19][9] = 4'hC;
    Number8[20][9] = 4'hC;
    Number8[21][9] = 4'hC;
    Number8[22][9] = 4'hF;
    Number8[23][9] = 4'hF;
    Number8[0][10] = 4'hF;
    Number8[1][10] = 4'hF;
    Number8[2][10] = 4'hC;
    Number8[3][10] = 4'hC;
    Number8[4][10] = 4'hC;
    Number8[5][10] = 4'hC;
    Number8[6][10] = 4'hC;
    Number8[7][10] = 4'hF;
    Number8[8][10] = 4'hF;
    Number8[9][10] = 4'hF;
    Number8[10][10] = 4'hF;
    Number8[11][10] = 4'hF;
    Number8[12][10] = 4'hF;
    Number8[13][10] = 4'hF;
    Number8[14][10] = 4'hF;
    Number8[15][10] = 4'hF;
    Number8[16][10] = 4'hF;
    Number8[17][10] = 4'hC;
    Number8[18][10] = 4'hC;
    Number8[19][10] = 4'hC;
    Number8[20][10] = 4'hC;
    Number8[21][10] = 4'hC;
    Number8[22][10] = 4'hF;
    Number8[23][10] = 4'hF;
    Number8[0][11] = 4'hF;
    Number8[1][11] = 4'hF;
    Number8[2][11] = 4'hC;
    Number8[3][11] = 4'hC;
    Number8[4][11] = 4'hC;
    Number8[5][11] = 4'hC;
    Number8[6][11] = 4'hC;
    Number8[7][11] = 4'hF;
    Number8[8][11] = 4'hF;
    Number8[9][11] = 4'hF;
    Number8[10][11] = 4'hF;
    Number8[11][11] = 4'hF;
    Number8[12][11] = 4'hF;
    Number8[13][11] = 4'hF;
    Number8[14][11] = 4'hF;
    Number8[15][11] = 4'hF;
    Number8[16][11] = 4'hF;
    Number8[17][11] = 4'hC;
    Number8[18][11] = 4'hC;
    Number8[19][11] = 4'hC;
    Number8[20][11] = 4'hC;
    Number8[21][11] = 4'hC;
    Number8[22][11] = 4'hF;
    Number8[23][11] = 4'hF;
    Number8[0][12] = 4'hF;
    Number8[1][12] = 4'hF;
    Number8[2][12] = 4'hC;
    Number8[3][12] = 4'hC;
    Number8[4][12] = 4'hC;
    Number8[5][12] = 4'hC;
    Number8[6][12] = 4'hC;
    Number8[7][12] = 4'hF;
    Number8[8][12] = 4'hF;
    Number8[9][12] = 4'hF;
    Number8[10][12] = 4'hF;
    Number8[11][12] = 4'hF;
    Number8[12][12] = 4'hF;
    Number8[13][12] = 4'hF;
    Number8[14][12] = 4'hF;
    Number8[15][12] = 4'hF;
    Number8[16][12] = 4'hF;
    Number8[17][12] = 4'hC;
    Number8[18][12] = 4'hC;
    Number8[19][12] = 4'hC;
    Number8[20][12] = 4'hC;
    Number8[21][12] = 4'hC;
    Number8[22][12] = 4'hF;
    Number8[23][12] = 4'hF;
    Number8[0][13] = 4'hF;
    Number8[1][13] = 4'hF;
    Number8[2][13] = 4'hF;
    Number8[3][13] = 4'hF;
    Number8[4][13] = 4'hF;
    Number8[5][13] = 4'hF;
    Number8[6][13] = 4'hF;
    Number8[7][13] = 4'hC;
    Number8[8][13] = 4'hC;
    Number8[9][13] = 4'hC;
    Number8[10][13] = 4'hC;
    Number8[11][13] = 4'hC;
    Number8[12][13] = 4'hC;
    Number8[13][13] = 4'hC;
    Number8[14][13] = 4'hC;
    Number8[15][13] = 4'hC;
    Number8[16][13] = 4'hC;
    Number8[17][13] = 4'hF;
    Number8[18][13] = 4'hF;
    Number8[19][13] = 4'hF;
    Number8[20][13] = 4'hF;
    Number8[21][13] = 4'hF;
    Number8[22][13] = 4'hF;
    Number8[23][13] = 4'hF;
    Number8[0][14] = 4'hF;
    Number8[1][14] = 4'hF;
    Number8[2][14] = 4'hF;
    Number8[3][14] = 4'hF;
    Number8[4][14] = 4'hF;
    Number8[5][14] = 4'hF;
    Number8[6][14] = 4'hF;
    Number8[7][14] = 4'hC;
    Number8[8][14] = 4'hC;
    Number8[9][14] = 4'hC;
    Number8[10][14] = 4'hC;
    Number8[11][14] = 4'hC;
    Number8[12][14] = 4'hC;
    Number8[13][14] = 4'hC;
    Number8[14][14] = 4'hC;
    Number8[15][14] = 4'hC;
    Number8[16][14] = 4'hC;
    Number8[17][14] = 4'hF;
    Number8[18][14] = 4'hF;
    Number8[19][14] = 4'hF;
    Number8[20][14] = 4'hF;
    Number8[21][14] = 4'hF;
    Number8[22][14] = 4'hF;
    Number8[23][14] = 4'hF;
    Number8[0][15] = 4'hF;
    Number8[1][15] = 4'hF;
    Number8[2][15] = 4'hF;
    Number8[3][15] = 4'hF;
    Number8[4][15] = 4'hF;
    Number8[5][15] = 4'hF;
    Number8[6][15] = 4'hF;
    Number8[7][15] = 4'hC;
    Number8[8][15] = 4'hC;
    Number8[9][15] = 4'hC;
    Number8[10][15] = 4'hC;
    Number8[11][15] = 4'hC;
    Number8[12][15] = 4'hC;
    Number8[13][15] = 4'hC;
    Number8[14][15] = 4'hC;
    Number8[15][15] = 4'hC;
    Number8[16][15] = 4'hC;
    Number8[17][15] = 4'hF;
    Number8[18][15] = 4'hF;
    Number8[19][15] = 4'hF;
    Number8[20][15] = 4'hF;
    Number8[21][15] = 4'hF;
    Number8[22][15] = 4'hF;
    Number8[23][15] = 4'hF;
    Number8[0][16] = 4'hF;
    Number8[1][16] = 4'hF;
    Number8[2][16] = 4'hF;
    Number8[3][16] = 4'hF;
    Number8[4][16] = 4'hF;
    Number8[5][16] = 4'hF;
    Number8[6][16] = 4'hF;
    Number8[7][16] = 4'hC;
    Number8[8][16] = 4'hC;
    Number8[9][16] = 4'hC;
    Number8[10][16] = 4'hC;
    Number8[11][16] = 4'hC;
    Number8[12][16] = 4'hC;
    Number8[13][16] = 4'hC;
    Number8[14][16] = 4'hC;
    Number8[15][16] = 4'hC;
    Number8[16][16] = 4'hC;
    Number8[17][16] = 4'hF;
    Number8[18][16] = 4'hF;
    Number8[19][16] = 4'hF;
    Number8[20][16] = 4'hF;
    Number8[21][16] = 4'hF;
    Number8[22][16] = 4'hF;
    Number8[23][16] = 4'hF;
    Number8[0][17] = 4'hF;
    Number8[1][17] = 4'hF;
    Number8[2][17] = 4'hF;
    Number8[3][17] = 4'hF;
    Number8[4][17] = 4'hF;
    Number8[5][17] = 4'hF;
    Number8[6][17] = 4'hF;
    Number8[7][17] = 4'hC;
    Number8[8][17] = 4'hC;
    Number8[9][17] = 4'hC;
    Number8[10][17] = 4'hC;
    Number8[11][17] = 4'hC;
    Number8[12][17] = 4'hC;
    Number8[13][17] = 4'hC;
    Number8[14][17] = 4'hC;
    Number8[15][17] = 4'hC;
    Number8[16][17] = 4'hC;
    Number8[17][17] = 4'hF;
    Number8[18][17] = 4'hF;
    Number8[19][17] = 4'hF;
    Number8[20][17] = 4'hF;
    Number8[21][17] = 4'hF;
    Number8[22][17] = 4'hF;
    Number8[23][17] = 4'hF;
    Number8[0][18] = 4'hF;
    Number8[1][18] = 4'hF;
    Number8[2][18] = 4'hC;
    Number8[3][18] = 4'hC;
    Number8[4][18] = 4'hC;
    Number8[5][18] = 4'hC;
    Number8[6][18] = 4'hC;
    Number8[7][18] = 4'hF;
    Number8[8][18] = 4'hF;
    Number8[9][18] = 4'hF;
    Number8[10][18] = 4'hF;
    Number8[11][18] = 4'hF;
    Number8[12][18] = 4'hF;
    Number8[13][18] = 4'hF;
    Number8[14][18] = 4'hF;
    Number8[15][18] = 4'hF;
    Number8[16][18] = 4'hF;
    Number8[17][18] = 4'hC;
    Number8[18][18] = 4'hC;
    Number8[19][18] = 4'hC;
    Number8[20][18] = 4'hC;
    Number8[21][18] = 4'hC;
    Number8[22][18] = 4'hF;
    Number8[23][18] = 4'hF;
    Number8[0][19] = 4'hF;
    Number8[1][19] = 4'hF;
    Number8[2][19] = 4'hC;
    Number8[3][19] = 4'hC;
    Number8[4][19] = 4'hC;
    Number8[5][19] = 4'hC;
    Number8[6][19] = 4'hC;
    Number8[7][19] = 4'hF;
    Number8[8][19] = 4'hF;
    Number8[9][19] = 4'hF;
    Number8[10][19] = 4'hF;
    Number8[11][19] = 4'hF;
    Number8[12][19] = 4'hF;
    Number8[13][19] = 4'hF;
    Number8[14][19] = 4'hF;
    Number8[15][19] = 4'hF;
    Number8[16][19] = 4'hF;
    Number8[17][19] = 4'hC;
    Number8[18][19] = 4'hC;
    Number8[19][19] = 4'hC;
    Number8[20][19] = 4'hC;
    Number8[21][19] = 4'hC;
    Number8[22][19] = 4'hF;
    Number8[23][19] = 4'hF;
    Number8[0][20] = 4'hF;
    Number8[1][20] = 4'hF;
    Number8[2][20] = 4'hC;
    Number8[3][20] = 4'hC;
    Number8[4][20] = 4'hC;
    Number8[5][20] = 4'hC;
    Number8[6][20] = 4'hC;
    Number8[7][20] = 4'hF;
    Number8[8][20] = 4'hF;
    Number8[9][20] = 4'hF;
    Number8[10][20] = 4'hF;
    Number8[11][20] = 4'hF;
    Number8[12][20] = 4'hF;
    Number8[13][20] = 4'hF;
    Number8[14][20] = 4'hF;
    Number8[15][20] = 4'hF;
    Number8[16][20] = 4'hF;
    Number8[17][20] = 4'hC;
    Number8[18][20] = 4'hC;
    Number8[19][20] = 4'hC;
    Number8[20][20] = 4'hC;
    Number8[21][20] = 4'hC;
    Number8[22][20] = 4'hF;
    Number8[23][20] = 4'hF;
    Number8[0][21] = 4'hF;
    Number8[1][21] = 4'hF;
    Number8[2][21] = 4'hC;
    Number8[3][21] = 4'hC;
    Number8[4][21] = 4'hC;
    Number8[5][21] = 4'hC;
    Number8[6][21] = 4'hC;
    Number8[7][21] = 4'hF;
    Number8[8][21] = 4'hF;
    Number8[9][21] = 4'hF;
    Number8[10][21] = 4'hF;
    Number8[11][21] = 4'hF;
    Number8[12][21] = 4'hF;
    Number8[13][21] = 4'hF;
    Number8[14][21] = 4'hF;
    Number8[15][21] = 4'hF;
    Number8[16][21] = 4'hF;
    Number8[17][21] = 4'hC;
    Number8[18][21] = 4'hC;
    Number8[19][21] = 4'hC;
    Number8[20][21] = 4'hC;
    Number8[21][21] = 4'hC;
    Number8[22][21] = 4'hF;
    Number8[23][21] = 4'hF;
    Number8[0][22] = 4'hF;
    Number8[1][22] = 4'hF;
    Number8[2][22] = 4'hC;
    Number8[3][22] = 4'hC;
    Number8[4][22] = 4'hC;
    Number8[5][22] = 4'hC;
    Number8[6][22] = 4'hC;
    Number8[7][22] = 4'hF;
    Number8[8][22] = 4'hF;
    Number8[9][22] = 4'hF;
    Number8[10][22] = 4'hF;
    Number8[11][22] = 4'hF;
    Number8[12][22] = 4'hF;
    Number8[13][22] = 4'hF;
    Number8[14][22] = 4'hF;
    Number8[15][22] = 4'hF;
    Number8[16][22] = 4'hF;
    Number8[17][22] = 4'hC;
    Number8[18][22] = 4'hC;
    Number8[19][22] = 4'hC;
    Number8[20][22] = 4'hC;
    Number8[21][22] = 4'hC;
    Number8[22][22] = 4'hF;
    Number8[23][22] = 4'hF;
    Number8[0][23] = 4'hF;
    Number8[1][23] = 4'hF;
    Number8[2][23] = 4'hF;
    Number8[3][23] = 4'hF;
    Number8[4][23] = 4'hF;
    Number8[5][23] = 4'hF;
    Number8[6][23] = 4'hF;
    Number8[7][23] = 4'hC;
    Number8[8][23] = 4'hC;
    Number8[9][23] = 4'hC;
    Number8[10][23] = 4'hC;
    Number8[11][23] = 4'hC;
    Number8[12][23] = 4'hC;
    Number8[13][23] = 4'hC;
    Number8[14][23] = 4'hC;
    Number8[15][23] = 4'hC;
    Number8[16][23] = 4'hC;
    Number8[17][23] = 4'hF;
    Number8[18][23] = 4'hF;
    Number8[19][23] = 4'hF;
    Number8[20][23] = 4'hF;
    Number8[21][23] = 4'hF;
    Number8[22][23] = 4'hF;
    Number8[23][23] = 4'hF;
    Number8[0][24] = 4'hF;
    Number8[1][24] = 4'hF;
    Number8[2][24] = 4'hF;
    Number8[3][24] = 4'hF;
    Number8[4][24] = 4'hF;
    Number8[5][24] = 4'hF;
    Number8[6][24] = 4'hF;
    Number8[7][24] = 4'hC;
    Number8[8][24] = 4'hC;
    Number8[9][24] = 4'hC;
    Number8[10][24] = 4'hC;
    Number8[11][24] = 4'hC;
    Number8[12][24] = 4'hC;
    Number8[13][24] = 4'hC;
    Number8[14][24] = 4'hC;
    Number8[15][24] = 4'hC;
    Number8[16][24] = 4'hC;
    Number8[17][24] = 4'hF;
    Number8[18][24] = 4'hF;
    Number8[19][24] = 4'hF;
    Number8[20][24] = 4'hF;
    Number8[21][24] = 4'hF;
    Number8[22][24] = 4'hF;
    Number8[23][24] = 4'hF;
    Number8[0][25] = 4'hF;
    Number8[1][25] = 4'hF;
    Number8[2][25] = 4'hF;
    Number8[3][25] = 4'hF;
    Number8[4][25] = 4'hF;
    Number8[5][25] = 4'hF;
    Number8[6][25] = 4'hF;
    Number8[7][25] = 4'hC;
    Number8[8][25] = 4'hC;
    Number8[9][25] = 4'hC;
    Number8[10][25] = 4'hC;
    Number8[11][25] = 4'hC;
    Number8[12][25] = 4'hC;
    Number8[13][25] = 4'hC;
    Number8[14][25] = 4'hC;
    Number8[15][25] = 4'hC;
    Number8[16][25] = 4'hC;
    Number8[17][25] = 4'hF;
    Number8[18][25] = 4'hF;
    Number8[19][25] = 4'hF;
    Number8[20][25] = 4'hF;
    Number8[21][25] = 4'hF;
    Number8[22][25] = 4'hF;
    Number8[23][25] = 4'hF;
    Number8[0][26] = 4'hF;
    Number8[1][26] = 4'hF;
    Number8[2][26] = 4'hF;
    Number8[3][26] = 4'hF;
    Number8[4][26] = 4'hF;
    Number8[5][26] = 4'hF;
    Number8[6][26] = 4'hF;
    Number8[7][26] = 4'hC;
    Number8[8][26] = 4'hC;
    Number8[9][26] = 4'hC;
    Number8[10][26] = 4'hC;
    Number8[11][26] = 4'hC;
    Number8[12][26] = 4'hC;
    Number8[13][26] = 4'hC;
    Number8[14][26] = 4'hC;
    Number8[15][26] = 4'hC;
    Number8[16][26] = 4'hC;
    Number8[17][26] = 4'hF;
    Number8[18][26] = 4'hF;
    Number8[19][26] = 4'hF;
    Number8[20][26] = 4'hF;
    Number8[21][26] = 4'hF;
    Number8[22][26] = 4'hF;
    Number8[23][26] = 4'hF;
    Number8[0][27] = 4'hF;
    Number8[1][27] = 4'hF;
    Number8[2][27] = 4'hF;
    Number8[3][27] = 4'hF;
    Number8[4][27] = 4'hF;
    Number8[5][27] = 4'hF;
    Number8[6][27] = 4'hF;
    Number8[7][27] = 4'hC;
    Number8[8][27] = 4'hC;
    Number8[9][27] = 4'hC;
    Number8[10][27] = 4'hC;
    Number8[11][27] = 4'hC;
    Number8[12][27] = 4'hC;
    Number8[13][27] = 4'hC;
    Number8[14][27] = 4'hC;
    Number8[15][27] = 4'hC;
    Number8[16][27] = 4'hC;
    Number8[17][27] = 4'hF;
    Number8[18][27] = 4'hF;
    Number8[19][27] = 4'hF;
    Number8[20][27] = 4'hF;
    Number8[21][27] = 4'hF;
    Number8[22][27] = 4'hF;
    Number8[23][27] = 4'hF;
    Number8[0][28] = 4'hF;
    Number8[1][28] = 4'hF;
    Number8[2][28] = 4'hF;
    Number8[3][28] = 4'hF;
    Number8[4][28] = 4'hF;
    Number8[5][28] = 4'hF;
    Number8[6][28] = 4'hF;
    Number8[7][28] = 4'hF;
    Number8[8][28] = 4'hF;
    Number8[9][28] = 4'hF;
    Number8[10][28] = 4'hF;
    Number8[11][28] = 4'hF;
    Number8[12][28] = 4'hF;
    Number8[13][28] = 4'hF;
    Number8[14][28] = 4'hF;
    Number8[15][28] = 4'hF;
    Number8[16][28] = 4'hF;
    Number8[17][28] = 4'hF;
    Number8[18][28] = 4'hF;
    Number8[19][28] = 4'hF;
    Number8[20][28] = 4'hF;
    Number8[21][28] = 4'hF;
    Number8[22][28] = 4'hF;
    Number8[23][28] = 4'hF;
    Number8[0][29] = 4'hF;
    Number8[1][29] = 4'hF;
    Number8[2][29] = 4'hF;
    Number8[3][29] = 4'hF;
    Number8[4][29] = 4'hF;
    Number8[5][29] = 4'hF;
    Number8[6][29] = 4'hF;
    Number8[7][29] = 4'hF;
    Number8[8][29] = 4'hF;
    Number8[9][29] = 4'hF;
    Number8[10][29] = 4'hF;
    Number8[11][29] = 4'hF;
    Number8[12][29] = 4'hF;
    Number8[13][29] = 4'hF;
    Number8[14][29] = 4'hF;
    Number8[15][29] = 4'hF;
    Number8[16][29] = 4'hF;
    Number8[17][29] = 4'hF;
    Number8[18][29] = 4'hF;
    Number8[19][29] = 4'hF;
    Number8[20][29] = 4'hF;
    Number8[21][29] = 4'hF;
    Number8[22][29] = 4'hF;
    Number8[23][29] = 4'hF;
 
//Number 9
    Number9[0][0] = 4'hF;
    Number9[1][0] = 4'hF;
    Number9[2][0] = 4'hF;
    Number9[3][0] = 4'hF;
    Number9[4][0] = 4'hF;
    Number9[5][0] = 4'hF;
    Number9[6][0] = 4'hF;
    Number9[7][0] = 4'hF;
    Number9[8][0] = 4'hF;
    Number9[9][0] = 4'hF;
    Number9[10][0] = 4'hF;
    Number9[11][0] = 4'hF;
    Number9[12][0] = 4'hF;
    Number9[13][0] = 4'hF;
    Number9[14][0] = 4'hF;
    Number9[15][0] = 4'hF;
    Number9[16][0] = 4'hF;
    Number9[17][0] = 4'hF;
    Number9[18][0] = 4'hF;
    Number9[19][0] = 4'hF;
    Number9[20][0] = 4'hF;
    Number9[21][0] = 4'hF;
    Number9[22][0] = 4'hF;
    Number9[23][0] = 4'hF;
    Number9[0][1] = 4'hF;
    Number9[1][1] = 4'hF;
    Number9[2][1] = 4'hF;
    Number9[3][1] = 4'hF;
    Number9[4][1] = 4'hF;
    Number9[5][1] = 4'hF;
    Number9[6][1] = 4'hF;
    Number9[7][1] = 4'hF;
    Number9[8][1] = 4'hF;
    Number9[9][1] = 4'hF;
    Number9[10][1] = 4'hF;
    Number9[11][1] = 4'hF;
    Number9[12][1] = 4'hF;
    Number9[13][1] = 4'hF;
    Number9[14][1] = 4'hF;
    Number9[15][1] = 4'hF;
    Number9[16][1] = 4'hF;
    Number9[17][1] = 4'hF;
    Number9[18][1] = 4'hF;
    Number9[19][1] = 4'hF;
    Number9[20][1] = 4'hF;
    Number9[21][1] = 4'hF;
    Number9[22][1] = 4'hF;
    Number9[23][1] = 4'hF;
    Number9[0][2] = 4'hF;
    Number9[1][2] = 4'hF;
    Number9[2][2] = 4'hF;
    Number9[3][2] = 4'hF;
    Number9[4][2] = 4'hF;
    Number9[5][2] = 4'hF;
    Number9[6][2] = 4'hF;
    Number9[7][2] = 4'hF;
    Number9[8][2] = 4'hF;
    Number9[9][2] = 4'hF;
    Number9[10][2] = 4'hF;
    Number9[11][2] = 4'hF;
    Number9[12][2] = 4'hF;
    Number9[13][2] = 4'hF;
    Number9[14][2] = 4'hF;
    Number9[15][2] = 4'hF;
    Number9[16][2] = 4'hF;
    Number9[17][2] = 4'hF;
    Number9[18][2] = 4'hF;
    Number9[19][2] = 4'hF;
    Number9[20][2] = 4'hF;
    Number9[21][2] = 4'hF;
    Number9[22][2] = 4'hF;
    Number9[23][2] = 4'hF;
    Number9[0][3] = 4'hF;
    Number9[1][3] = 4'hF;
    Number9[2][3] = 4'hF;
    Number9[3][3] = 4'hF;
    Number9[4][3] = 4'hF;
    Number9[5][3] = 4'hF;
    Number9[6][3] = 4'hF;
    Number9[7][3] = 4'hC;
    Number9[8][3] = 4'hC;
    Number9[9][3] = 4'hC;
    Number9[10][3] = 4'hC;
    Number9[11][3] = 4'hC;
    Number9[12][3] = 4'hC;
    Number9[13][3] = 4'hC;
    Number9[14][3] = 4'hC;
    Number9[15][3] = 4'hC;
    Number9[16][3] = 4'hC;
    Number9[17][3] = 4'hF;
    Number9[18][3] = 4'hF;
    Number9[19][3] = 4'hF;
    Number9[20][3] = 4'hF;
    Number9[21][3] = 4'hF;
    Number9[22][3] = 4'hF;
    Number9[23][3] = 4'hF;
    Number9[0][4] = 4'hF;
    Number9[1][4] = 4'hF;
    Number9[2][4] = 4'hF;
    Number9[3][4] = 4'hF;
    Number9[4][4] = 4'hF;
    Number9[5][4] = 4'hF;
    Number9[6][4] = 4'hF;
    Number9[7][4] = 4'hC;
    Number9[8][4] = 4'hC;
    Number9[9][4] = 4'hC;
    Number9[10][4] = 4'hC;
    Number9[11][4] = 4'hC;
    Number9[12][4] = 4'hC;
    Number9[13][4] = 4'hC;
    Number9[14][4] = 4'hC;
    Number9[15][4] = 4'hC;
    Number9[16][4] = 4'hC;
    Number9[17][4] = 4'hF;
    Number9[18][4] = 4'hF;
    Number9[19][4] = 4'hF;
    Number9[20][4] = 4'hF;
    Number9[21][4] = 4'hF;
    Number9[22][4] = 4'hF;
    Number9[23][4] = 4'hF;
    Number9[0][5] = 4'hF;
    Number9[1][5] = 4'hF;
    Number9[2][5] = 4'hF;
    Number9[3][5] = 4'hF;
    Number9[4][5] = 4'hF;
    Number9[5][5] = 4'hF;
    Number9[6][5] = 4'hF;
    Number9[7][5] = 4'hC;
    Number9[8][5] = 4'hC;
    Number9[9][5] = 4'hC;
    Number9[10][5] = 4'hC;
    Number9[11][5] = 4'hC;
    Number9[12][5] = 4'hC;
    Number9[13][5] = 4'hC;
    Number9[14][5] = 4'hC;
    Number9[15][5] = 4'hC;
    Number9[16][5] = 4'hC;
    Number9[17][5] = 4'hF;
    Number9[18][5] = 4'hF;
    Number9[19][5] = 4'hF;
    Number9[20][5] = 4'hF;
    Number9[21][5] = 4'hF;
    Number9[22][5] = 4'hF;
    Number9[23][5] = 4'hF;
    Number9[0][6] = 4'hF;
    Number9[1][6] = 4'hF;
    Number9[2][6] = 4'hF;
    Number9[3][6] = 4'hF;
    Number9[4][6] = 4'hF;
    Number9[5][6] = 4'hF;
    Number9[6][6] = 4'hF;
    Number9[7][6] = 4'hC;
    Number9[8][6] = 4'hC;
    Number9[9][6] = 4'hC;
    Number9[10][6] = 4'hC;
    Number9[11][6] = 4'hC;
    Number9[12][6] = 4'hC;
    Number9[13][6] = 4'hC;
    Number9[14][6] = 4'hC;
    Number9[15][6] = 4'hC;
    Number9[16][6] = 4'hC;
    Number9[17][6] = 4'hF;
    Number9[18][6] = 4'hF;
    Number9[19][6] = 4'hF;
    Number9[20][6] = 4'hF;
    Number9[21][6] = 4'hF;
    Number9[22][6] = 4'hF;
    Number9[23][6] = 4'hF;
    Number9[0][7] = 4'hF;
    Number9[1][7] = 4'hF;
    Number9[2][7] = 4'hF;
    Number9[3][7] = 4'hF;
    Number9[4][7] = 4'hF;
    Number9[5][7] = 4'hF;
    Number9[6][7] = 4'hF;
    Number9[7][7] = 4'hC;
    Number9[8][7] = 4'hC;
    Number9[9][7] = 4'hC;
    Number9[10][7] = 4'hC;
    Number9[11][7] = 4'hC;
    Number9[12][7] = 4'hC;
    Number9[13][7] = 4'hC;
    Number9[14][7] = 4'hC;
    Number9[15][7] = 4'hC;
    Number9[16][7] = 4'hC;
    Number9[17][7] = 4'hF;
    Number9[18][7] = 4'hF;
    Number9[19][7] = 4'hF;
    Number9[20][7] = 4'hF;
    Number9[21][7] = 4'hF;
    Number9[22][7] = 4'hF;
    Number9[23][7] = 4'hF;
    Number9[0][8] = 4'hF;
    Number9[1][8] = 4'hF;
    Number9[2][8] = 4'hC;
    Number9[3][8] = 4'hC;
    Number9[4][8] = 4'hC;
    Number9[5][8] = 4'hC;
    Number9[6][8] = 4'hC;
    Number9[7][8] = 4'hF;
    Number9[8][8] = 4'hF;
    Number9[9][8] = 4'hF;
    Number9[10][8] = 4'hF;
    Number9[11][8] = 4'hF;
    Number9[12][8] = 4'hF;
    Number9[13][8] = 4'hF;
    Number9[14][8] = 4'hF;
    Number9[15][8] = 4'hF;
    Number9[16][8] = 4'hF;
    Number9[17][8] = 4'hC;
    Number9[18][8] = 4'hC;
    Number9[19][8] = 4'hC;
    Number9[20][8] = 4'hC;
    Number9[21][8] = 4'hC;
    Number9[22][8] = 4'hF;
    Number9[23][8] = 4'hF;
    Number9[0][9] = 4'hF;
    Number9[1][9] = 4'hF;
    Number9[2][9] = 4'hC;
    Number9[3][9] = 4'hC;
    Number9[4][9] = 4'hC;
    Number9[5][9] = 4'hC;
    Number9[6][9] = 4'hC;
    Number9[7][9] = 4'hF;
    Number9[8][9] = 4'hF;
    Number9[9][9] = 4'hF;
    Number9[10][9] = 4'hF;
    Number9[11][9] = 4'hF;
    Number9[12][9] = 4'hF;
    Number9[13][9] = 4'hF;
    Number9[14][9] = 4'hF;
    Number9[15][9] = 4'hF;
    Number9[16][9] = 4'hF;
    Number9[17][9] = 4'hC;
    Number9[18][9] = 4'hC;
    Number9[19][9] = 4'hC;
    Number9[20][9] = 4'hC;
    Number9[21][9] = 4'hC;
    Number9[22][9] = 4'hF;
    Number9[23][9] = 4'hF;
    Number9[0][10] = 4'hF;
    Number9[1][10] = 4'hF;
    Number9[2][10] = 4'hC;
    Number9[3][10] = 4'hC;
    Number9[4][10] = 4'hC;
    Number9[5][10] = 4'hC;
    Number9[6][10] = 4'hC;
    Number9[7][10] = 4'hF;
    Number9[8][10] = 4'hF;
    Number9[9][10] = 4'hF;
    Number9[10][10] = 4'hF;
    Number9[11][10] = 4'hF;
    Number9[12][10] = 4'hF;
    Number9[13][10] = 4'hF;
    Number9[14][10] = 4'hF;
    Number9[15][10] = 4'hF;
    Number9[16][10] = 4'hF;
    Number9[17][10] = 4'hC;
    Number9[18][10] = 4'hC;
    Number9[19][10] = 4'hC;
    Number9[20][10] = 4'hC;
    Number9[21][10] = 4'hC;
    Number9[22][10] = 4'hF;
    Number9[23][10] = 4'hF;
    Number9[0][11] = 4'hF;
    Number9[1][11] = 4'hF;
    Number9[2][11] = 4'hC;
    Number9[3][11] = 4'hC;
    Number9[4][11] = 4'hC;
    Number9[5][11] = 4'hC;
    Number9[6][11] = 4'hC;
    Number9[7][11] = 4'hF;
    Number9[8][11] = 4'hF;
    Number9[9][11] = 4'hF;
    Number9[10][11] = 4'hF;
    Number9[11][11] = 4'hF;
    Number9[12][11] = 4'hF;
    Number9[13][11] = 4'hF;
    Number9[14][11] = 4'hF;
    Number9[15][11] = 4'hF;
    Number9[16][11] = 4'hF;
    Number9[17][11] = 4'hC;
    Number9[18][11] = 4'hC;
    Number9[19][11] = 4'hC;
    Number9[20][11] = 4'hC;
    Number9[21][11] = 4'hC;
    Number9[22][11] = 4'hF;
    Number9[23][11] = 4'hF;
    Number9[0][12] = 4'hF;
    Number9[1][12] = 4'hF;
    Number9[2][12] = 4'hC;
    Number9[3][12] = 4'hC;
    Number9[4][12] = 4'hC;
    Number9[5][12] = 4'hC;
    Number9[6][12] = 4'hC;
    Number9[7][12] = 4'hF;
    Number9[8][12] = 4'hF;
    Number9[9][12] = 4'hF;
    Number9[10][12] = 4'hF;
    Number9[11][12] = 4'hF;
    Number9[12][12] = 4'hF;
    Number9[13][12] = 4'hF;
    Number9[14][12] = 4'hF;
    Number9[15][12] = 4'hF;
    Number9[16][12] = 4'hF;
    Number9[17][12] = 4'hC;
    Number9[18][12] = 4'hC;
    Number9[19][12] = 4'hC;
    Number9[20][12] = 4'hC;
    Number9[21][12] = 4'hC;
    Number9[22][12] = 4'hF;
    Number9[23][12] = 4'hF;
    Number9[0][13] = 4'hF;
    Number9[1][13] = 4'hF;
    Number9[2][13] = 4'hF;
    Number9[3][13] = 4'hF;
    Number9[4][13] = 4'hF;
    Number9[5][13] = 4'hF;
    Number9[6][13] = 4'hF;
    Number9[7][13] = 4'hC;
    Number9[8][13] = 4'hC;
    Number9[9][13] = 4'hC;
    Number9[10][13] = 4'hC;
    Number9[11][13] = 4'hC;
    Number9[12][13] = 4'hC;
    Number9[13][13] = 4'hC;
    Number9[14][13] = 4'hC;
    Number9[15][13] = 4'hC;
    Number9[16][13] = 4'hC;
    Number9[17][13] = 4'hC;
    Number9[18][13] = 4'hC;
    Number9[19][13] = 4'hC;
    Number9[20][13] = 4'hC;
    Number9[21][13] = 4'hC;
    Number9[22][13] = 4'hF;
    Number9[23][13] = 4'hF;
    Number9[0][14] = 4'hF;
    Number9[1][14] = 4'hF;
    Number9[2][14] = 4'hF;
    Number9[3][14] = 4'hF;
    Number9[4][14] = 4'hF;
    Number9[5][14] = 4'hF;
    Number9[6][14] = 4'hF;
    Number9[7][14] = 4'hC;
    Number9[8][14] = 4'hC;
    Number9[9][14] = 4'hC;
    Number9[10][14] = 4'hC;
    Number9[11][14] = 4'hC;
    Number9[12][14] = 4'hC;
    Number9[13][14] = 4'hC;
    Number9[14][14] = 4'hC;
    Number9[15][14] = 4'hC;
    Number9[16][14] = 4'hC;
    Number9[17][14] = 4'hC;
    Number9[18][14] = 4'hC;
    Number9[19][14] = 4'hC;
    Number9[20][14] = 4'hC;
    Number9[21][14] = 4'hC;
    Number9[22][14] = 4'hF;
    Number9[23][14] = 4'hF;
    Number9[0][15] = 4'hF;
    Number9[1][15] = 4'hF;
    Number9[2][15] = 4'hF;
    Number9[3][15] = 4'hF;
    Number9[4][15] = 4'hF;
    Number9[5][15] = 4'hF;
    Number9[6][15] = 4'hF;
    Number9[7][15] = 4'hC;
    Number9[8][15] = 4'hC;
    Number9[9][15] = 4'hC;
    Number9[10][15] = 4'hC;
    Number9[11][15] = 4'hC;
    Number9[12][15] = 4'hC;
    Number9[13][15] = 4'hC;
    Number9[14][15] = 4'hC;
    Number9[15][15] = 4'hC;
    Number9[16][15] = 4'hC;
    Number9[17][15] = 4'hC;
    Number9[18][15] = 4'hC;
    Number9[19][15] = 4'hC;
    Number9[20][15] = 4'hC;
    Number9[21][15] = 4'hC;
    Number9[22][15] = 4'hF;
    Number9[23][15] = 4'hF;
    Number9[0][16] = 4'hF;
    Number9[1][16] = 4'hF;
    Number9[2][16] = 4'hF;
    Number9[3][16] = 4'hF;
    Number9[4][16] = 4'hF;
    Number9[5][16] = 4'hF;
    Number9[6][16] = 4'hF;
    Number9[7][16] = 4'hC;
    Number9[8][16] = 4'hC;
    Number9[9][16] = 4'hC;
    Number9[10][16] = 4'hC;
    Number9[11][16] = 4'hC;
    Number9[12][16] = 4'hC;
    Number9[13][16] = 4'hC;
    Number9[14][16] = 4'hC;
    Number9[15][16] = 4'hC;
    Number9[16][16] = 4'hC;
    Number9[17][16] = 4'hC;
    Number9[18][16] = 4'hC;
    Number9[19][16] = 4'hC;
    Number9[20][16] = 4'hC;
    Number9[21][16] = 4'hC;
    Number9[22][16] = 4'hF;
    Number9[23][16] = 4'hF;
    Number9[0][17] = 4'hF;
    Number9[1][17] = 4'hF;
    Number9[2][17] = 4'hF;
    Number9[3][17] = 4'hF;
    Number9[4][17] = 4'hF;
    Number9[5][17] = 4'hF;
    Number9[6][17] = 4'hF;
    Number9[7][17] = 4'hC;
    Number9[8][17] = 4'hC;
    Number9[9][17] = 4'hC;
    Number9[10][17] = 4'hC;
    Number9[11][17] = 4'hC;
    Number9[12][17] = 4'hC;
    Number9[13][17] = 4'hC;
    Number9[14][17] = 4'hC;
    Number9[15][17] = 4'hC;
    Number9[16][17] = 4'hC;
    Number9[17][17] = 4'hC;
    Number9[18][17] = 4'hC;
    Number9[19][17] = 4'hC;
    Number9[20][17] = 4'hC;
    Number9[21][17] = 4'hC;
    Number9[22][17] = 4'hF;
    Number9[23][17] = 4'hF;
    Number9[0][18] = 4'hF;
    Number9[1][18] = 4'hF;
    Number9[2][18] = 4'hF;
    Number9[3][18] = 4'hF;
    Number9[4][18] = 4'hF;
    Number9[5][18] = 4'hF;
    Number9[6][18] = 4'hF;
    Number9[7][18] = 4'hF;
    Number9[8][18] = 4'hF;
    Number9[9][18] = 4'hF;
    Number9[10][18] = 4'hF;
    Number9[11][18] = 4'hF;
    Number9[12][18] = 4'hF;
    Number9[13][18] = 4'hF;
    Number9[14][18] = 4'hF;
    Number9[15][18] = 4'hF;
    Number9[16][18] = 4'hF;
    Number9[17][18] = 4'hC;
    Number9[18][18] = 4'hC;
    Number9[19][18] = 4'hC;
    Number9[20][18] = 4'hC;
    Number9[21][18] = 4'hC;
    Number9[22][18] = 4'hF;
    Number9[23][18] = 4'hF;
    Number9[0][19] = 4'hF;
    Number9[1][19] = 4'hF;
    Number9[2][19] = 4'hF;
    Number9[3][19] = 4'hF;
    Number9[4][19] = 4'hF;
    Number9[5][19] = 4'hF;
    Number9[6][19] = 4'hF;
    Number9[7][19] = 4'hF;
    Number9[8][19] = 4'hF;
    Number9[9][19] = 4'hF;
    Number9[10][19] = 4'hF;
    Number9[11][19] = 4'hF;
    Number9[12][19] = 4'hF;
    Number9[13][19] = 4'hF;
    Number9[14][19] = 4'hF;
    Number9[15][19] = 4'hF;
    Number9[16][19] = 4'hF;
    Number9[17][19] = 4'hC;
    Number9[18][19] = 4'hC;
    Number9[19][19] = 4'hC;
    Number9[20][19] = 4'hC;
    Number9[21][19] = 4'hC;
    Number9[22][19] = 4'hF;
    Number9[23][19] = 4'hF;
    Number9[0][20] = 4'hF;
    Number9[1][20] = 4'hF;
    Number9[2][20] = 4'hF;
    Number9[3][20] = 4'hF;
    Number9[4][20] = 4'hF;
    Number9[5][20] = 4'hF;
    Number9[6][20] = 4'hF;
    Number9[7][20] = 4'hF;
    Number9[8][20] = 4'hF;
    Number9[9][20] = 4'hF;
    Number9[10][20] = 4'hF;
    Number9[11][20] = 4'hF;
    Number9[12][20] = 4'hF;
    Number9[13][20] = 4'hF;
    Number9[14][20] = 4'hF;
    Number9[15][20] = 4'hF;
    Number9[16][20] = 4'hF;
    Number9[17][20] = 4'hC;
    Number9[18][20] = 4'hC;
    Number9[19][20] = 4'hC;
    Number9[20][20] = 4'hC;
    Number9[21][20] = 4'hC;
    Number9[22][20] = 4'hF;
    Number9[23][20] = 4'hF;
    Number9[0][21] = 4'hF;
    Number9[1][21] = 4'hF;
    Number9[2][21] = 4'hF;
    Number9[3][21] = 4'hF;
    Number9[4][21] = 4'hF;
    Number9[5][21] = 4'hF;
    Number9[6][21] = 4'hF;
    Number9[7][21] = 4'hF;
    Number9[8][21] = 4'hF;
    Number9[9][21] = 4'hF;
    Number9[10][21] = 4'hF;
    Number9[11][21] = 4'hF;
    Number9[12][21] = 4'hF;
    Number9[13][21] = 4'hF;
    Number9[14][21] = 4'hF;
    Number9[15][21] = 4'hF;
    Number9[16][21] = 4'hF;
    Number9[17][21] = 4'hC;
    Number9[18][21] = 4'hC;
    Number9[19][21] = 4'hC;
    Number9[20][21] = 4'hC;
    Number9[21][21] = 4'hC;
    Number9[22][21] = 4'hF;
    Number9[23][21] = 4'hF;
    Number9[0][22] = 4'hF;
    Number9[1][22] = 4'hF;
    Number9[2][22] = 4'hF;
    Number9[3][22] = 4'hF;
    Number9[4][22] = 4'hF;
    Number9[5][22] = 4'hF;
    Number9[6][22] = 4'hF;
    Number9[7][22] = 4'hF;
    Number9[8][22] = 4'hF;
    Number9[9][22] = 4'hF;
    Number9[10][22] = 4'hF;
    Number9[11][22] = 4'hF;
    Number9[12][22] = 4'hF;
    Number9[13][22] = 4'hF;
    Number9[14][22] = 4'hF;
    Number9[15][22] = 4'hF;
    Number9[16][22] = 4'hF;
    Number9[17][22] = 4'hC;
    Number9[18][22] = 4'hC;
    Number9[19][22] = 4'hC;
    Number9[20][22] = 4'hC;
    Number9[21][22] = 4'hC;
    Number9[22][22] = 4'hF;
    Number9[23][22] = 4'hF;
    Number9[0][23] = 4'hF;
    Number9[1][23] = 4'hF;
    Number9[2][23] = 4'hF;
    Number9[3][23] = 4'hF;
    Number9[4][23] = 4'hF;
    Number9[5][23] = 4'hF;
    Number9[6][23] = 4'hF;
    Number9[7][23] = 4'hC;
    Number9[8][23] = 4'hC;
    Number9[9][23] = 4'hC;
    Number9[10][23] = 4'hC;
    Number9[11][23] = 4'hC;
    Number9[12][23] = 4'hC;
    Number9[13][23] = 4'hC;
    Number9[14][23] = 4'hC;
    Number9[15][23] = 4'hC;
    Number9[16][23] = 4'hC;
    Number9[17][23] = 4'hF;
    Number9[18][23] = 4'hF;
    Number9[19][23] = 4'hF;
    Number9[20][23] = 4'hF;
    Number9[21][23] = 4'hF;
    Number9[22][23] = 4'hF;
    Number9[23][23] = 4'hF;
    Number9[0][24] = 4'hF;
    Number9[1][24] = 4'hF;
    Number9[2][24] = 4'hF;
    Number9[3][24] = 4'hF;
    Number9[4][24] = 4'hF;
    Number9[5][24] = 4'hF;
    Number9[6][24] = 4'hF;
    Number9[7][24] = 4'hC;
    Number9[8][24] = 4'hC;
    Number9[9][24] = 4'hC;
    Number9[10][24] = 4'hC;
    Number9[11][24] = 4'hC;
    Number9[12][24] = 4'hC;
    Number9[13][24] = 4'hC;
    Number9[14][24] = 4'hC;
    Number9[15][24] = 4'hC;
    Number9[16][24] = 4'hC;
    Number9[17][24] = 4'hF;
    Number9[18][24] = 4'hF;
    Number9[19][24] = 4'hF;
    Number9[20][24] = 4'hF;
    Number9[21][24] = 4'hF;
    Number9[22][24] = 4'hF;
    Number9[23][24] = 4'hF;
    Number9[0][25] = 4'hF;
    Number9[1][25] = 4'hF;
    Number9[2][25] = 4'hF;
    Number9[3][25] = 4'hF;
    Number9[4][25] = 4'hF;
    Number9[5][25] = 4'hF;
    Number9[6][25] = 4'hF;
    Number9[7][25] = 4'hC;
    Number9[8][25] = 4'hC;
    Number9[9][25] = 4'hC;
    Number9[10][25] = 4'hC;
    Number9[11][25] = 4'hC;
    Number9[12][25] = 4'hC;
    Number9[13][25] = 4'hC;
    Number9[14][25] = 4'hC;
    Number9[15][25] = 4'hC;
    Number9[16][25] = 4'hC;
    Number9[17][25] = 4'hF;
    Number9[18][25] = 4'hF;
    Number9[19][25] = 4'hF;
    Number9[20][25] = 4'hF;
    Number9[21][25] = 4'hF;
    Number9[22][25] = 4'hF;
    Number9[23][25] = 4'hF;
    Number9[0][26] = 4'hF;
    Number9[1][26] = 4'hF;
    Number9[2][26] = 4'hF;
    Number9[3][26] = 4'hF;
    Number9[4][26] = 4'hF;
    Number9[5][26] = 4'hF;
    Number9[6][26] = 4'hF;
    Number9[7][26] = 4'hC;
    Number9[8][26] = 4'hC;
    Number9[9][26] = 4'hC;
    Number9[10][26] = 4'hC;
    Number9[11][26] = 4'hC;
    Number9[12][26] = 4'hC;
    Number9[13][26] = 4'hC;
    Number9[14][26] = 4'hC;
    Number9[15][26] = 4'hC;
    Number9[16][26] = 4'hC;
    Number9[17][26] = 4'hF;
    Number9[18][26] = 4'hF;
    Number9[19][26] = 4'hF;
    Number9[20][26] = 4'hF;
    Number9[21][26] = 4'hF;
    Number9[22][26] = 4'hF;
    Number9[23][26] = 4'hF;
    Number9[0][27] = 4'hF;
    Number9[1][27] = 4'hF;
    Number9[2][27] = 4'hF;
    Number9[3][27] = 4'hF;
    Number9[4][27] = 4'hF;
    Number9[5][27] = 4'hF;
    Number9[6][27] = 4'hF;
    Number9[7][27] = 4'hC;
    Number9[8][27] = 4'hC;
    Number9[9][27] = 4'hC;
    Number9[10][27] = 4'hC;
    Number9[11][27] = 4'hC;
    Number9[12][27] = 4'hC;
    Number9[13][27] = 4'hC;
    Number9[14][27] = 4'hC;
    Number9[15][27] = 4'hC;
    Number9[16][27] = 4'hC;
    Number9[17][27] = 4'hF;
    Number9[18][27] = 4'hF;
    Number9[19][27] = 4'hF;
    Number9[20][27] = 4'hF;
    Number9[21][27] = 4'hF;
    Number9[22][27] = 4'hF;
    Number9[23][27] = 4'hF;
    Number9[0][28] = 4'hF;
    Number9[1][28] = 4'hF;
    Number9[2][28] = 4'hF;
    Number9[3][28] = 4'hF;
    Number9[4][28] = 4'hF;
    Number9[5][28] = 4'hF;
    Number9[6][28] = 4'hF;
    Number9[7][28] = 4'hF;
    Number9[8][28] = 4'hF;
    Number9[9][28] = 4'hF;
    Number9[10][28] = 4'hF;
    Number9[11][28] = 4'hF;
    Number9[12][28] = 4'hF;
    Number9[13][28] = 4'hF;
    Number9[14][28] = 4'hF;
    Number9[15][28] = 4'hF;
    Number9[16][28] = 4'hF;
    Number9[17][28] = 4'hF;
    Number9[18][28] = 4'hF;
    Number9[19][28] = 4'hF;
    Number9[20][28] = 4'hF;
    Number9[21][28] = 4'hF;
    Number9[22][28] = 4'hF;
    Number9[23][28] = 4'hF;
    Number9[0][29] = 4'hF;
    Number9[1][29] = 4'hF;
    Number9[2][29] = 4'hF;
    Number9[3][29] = 4'hF;
    Number9[4][29] = 4'hF;
    Number9[5][29] = 4'hF;
    Number9[6][29] = 4'hF;
    Number9[7][29] = 4'hF;
    Number9[8][29] = 4'hF;
    Number9[9][29] = 4'hF;
    Number9[10][29] = 4'hF;
    Number9[11][29] = 4'hF;
    Number9[12][29] = 4'hF;
    Number9[13][29] = 4'hF;
    Number9[14][29] = 4'hF;
    Number9[15][29] = 4'hF;
    Number9[16][29] = 4'hF;
    Number9[17][29] = 4'hF;
    Number9[18][29] = 4'hF;
    Number9[19][29] = 4'hF;
    Number9[20][29] = 4'hF;
    Number9[21][29] = 4'hF;
    Number9[22][29] = 4'hF;
    Number9[23][29] = 4'hF;

// Storing information about the Article images

// Score article 
    S_A[0][0] = 4'hF;
    S_A[1][0] = 4'hF;
    S_A[2][0] = 4'hF;
    S_A[3][0] = 4'hF;
    S_A[4][0] = 4'hF;
    S_A[5][0] = 4'hF;
    S_A[6][0] = 4'hF;
    S_A[7][0] = 4'hF;
    S_A[8][0] = 4'hF;
    S_A[9][0] = 4'hF;
    S_A[10][0] = 4'hF;
    S_A[11][0] = 4'hF;
    S_A[12][0] = 4'hF;
    S_A[13][0] = 4'hF;
    S_A[14][0] = 4'hF;
    S_A[15][0] = 4'hF;
    S_A[16][0] = 4'hF;
    S_A[17][0] = 4'hF;
    S_A[18][0] = 4'hF;
    S_A[19][0] = 4'hF;
    S_A[20][0] = 4'hF;
    S_A[21][0] = 4'hF;
    S_A[22][0] = 4'hF;
    S_A[23][0] = 4'hF;
    S_A[24][0] = 4'hF;
    S_A[25][0] = 4'hF;
    S_A[26][0] = 4'hF;
    S_A[27][0] = 4'hF;
    S_A[28][0] = 4'hF;
    S_A[29][0] = 4'hF;
    S_A[30][0] = 4'hF;
    S_A[31][0] = 4'hF;
    S_A[32][0] = 4'hF;
    S_A[33][0] = 4'hF;
    S_A[34][0] = 4'hF;
    S_A[35][0] = 4'hF;
    S_A[36][0] = 4'hF;
    S_A[37][0] = 4'hF;
    S_A[38][0] = 4'hF;
    S_A[39][0] = 4'hF;
    S_A[40][0] = 4'hF;
    S_A[41][0] = 4'hF;
    S_A[42][0] = 4'hF;
    S_A[43][0] = 4'hF;
    S_A[44][0] = 4'hF;
    S_A[45][0] = 4'hF;
    S_A[46][0] = 4'hF;
    S_A[47][0] = 4'hF;
    S_A[48][0] = 4'hF;
    S_A[49][0] = 4'hF;
    S_A[50][0] = 4'hF;
    S_A[51][0] = 4'hF;
    S_A[52][0] = 4'hF;
    S_A[53][0] = 4'hF;
    S_A[54][0] = 4'hF;
    S_A[55][0] = 4'hF;
    S_A[56][0] = 4'hF;
    S_A[57][0] = 4'hF;
    S_A[58][0] = 4'hF;
    S_A[59][0] = 4'hF;
    S_A[60][0] = 4'hF;
    S_A[61][0] = 4'hF;
    S_A[62][0] = 4'hF;
    S_A[63][0] = 4'hF;
    S_A[64][0] = 4'hF;
    S_A[65][0] = 4'hF;
    S_A[66][0] = 4'hF;
    S_A[67][0] = 4'hF;
    S_A[68][0] = 4'hF;
    S_A[69][0] = 4'hF;
    S_A[70][0] = 4'hF;
    S_A[71][0] = 4'hF;
    S_A[72][0] = 4'hF;
    S_A[73][0] = 4'hF;
    S_A[74][0] = 4'hF;
    S_A[75][0] = 4'hF;
    S_A[76][0] = 4'hF;
    S_A[77][0] = 4'hF;
    S_A[78][0] = 4'hF;
    S_A[79][0] = 4'hF;
    S_A[80][0] = 4'hF;
    S_A[81][0] = 4'hF;
    S_A[82][0] = 4'hF;
    S_A[83][0] = 4'hF;
    S_A[84][0] = 4'hF;
    S_A[85][0] = 4'hF;
    S_A[86][0] = 4'hF;
    S_A[87][0] = 4'hF;
    S_A[88][0] = 4'hF;
    S_A[89][0] = 4'hF;
    S_A[90][0] = 4'hF;
    S_A[91][0] = 4'hF;
    S_A[92][0] = 4'hF;
    S_A[93][0] = 4'hF;
    S_A[94][0] = 4'hF;
    S_A[95][0] = 4'hF;
    S_A[96][0] = 4'hF;
    S_A[97][0] = 4'hF;
    S_A[98][0] = 4'hF;
    S_A[99][0] = 4'hF;
    S_A[100][0] = 4'hF;
    S_A[101][0] = 4'hF;
    S_A[102][0] = 4'hF;
    S_A[103][0] = 4'hF;
    S_A[104][0] = 4'hF;
    S_A[105][0] = 4'hF;
    S_A[106][0] = 4'hF;
    S_A[107][0] = 4'hF;
    S_A[108][0] = 4'hF;
    S_A[109][0] = 4'hF;
    S_A[110][0] = 4'hF;
    S_A[111][0] = 4'hF;
    S_A[112][0] = 4'hF;
    S_A[113][0] = 4'hF;
    S_A[114][0] = 4'hF;
    S_A[0][1] = 4'hF;
    S_A[1][1] = 4'hF;
    S_A[2][1] = 4'hF;
    S_A[3][1] = 4'hF;
    S_A[4][1] = 4'hF;
    S_A[5][1] = 4'hF;
    S_A[6][1] = 4'hF;
    S_A[7][1] = 4'hF;
    S_A[8][1] = 4'hF;
    S_A[9][1] = 4'hF;
    S_A[10][1] = 4'hF;
    S_A[11][1] = 4'hF;
    S_A[12][1] = 4'hF;
    S_A[13][1] = 4'hF;
    S_A[14][1] = 4'hF;
    S_A[15][1] = 4'hF;
    S_A[16][1] = 4'hF;
    S_A[17][1] = 4'hF;
    S_A[18][1] = 4'hF;
    S_A[19][1] = 4'hF;
    S_A[20][1] = 4'hF;
    S_A[21][1] = 4'hF;
    S_A[22][1] = 4'hF;
    S_A[23][1] = 4'hF;
    S_A[24][1] = 4'hF;
    S_A[25][1] = 4'hF;
    S_A[26][1] = 4'hF;
    S_A[27][1] = 4'hF;
    S_A[28][1] = 4'hF;
    S_A[29][1] = 4'hF;
    S_A[30][1] = 4'hF;
    S_A[31][1] = 4'hF;
    S_A[32][1] = 4'hF;
    S_A[33][1] = 4'hF;
    S_A[34][1] = 4'hF;
    S_A[35][1] = 4'hF;
    S_A[36][1] = 4'hF;
    S_A[37][1] = 4'hF;
    S_A[38][1] = 4'hF;
    S_A[39][1] = 4'hF;
    S_A[40][1] = 4'hF;
    S_A[41][1] = 4'hF;
    S_A[42][1] = 4'hF;
    S_A[43][1] = 4'hF;
    S_A[44][1] = 4'hF;
    S_A[45][1] = 4'hF;
    S_A[46][1] = 4'hF;
    S_A[47][1] = 4'hF;
    S_A[48][1] = 4'hF;
    S_A[49][1] = 4'hF;
    S_A[50][1] = 4'hF;
    S_A[51][1] = 4'hF;
    S_A[52][1] = 4'hF;
    S_A[53][1] = 4'hF;
    S_A[54][1] = 4'hF;
    S_A[55][1] = 4'hF;
    S_A[56][1] = 4'hF;
    S_A[57][1] = 4'hF;
    S_A[58][1] = 4'hF;
    S_A[59][1] = 4'hF;
    S_A[60][1] = 4'hF;
    S_A[61][1] = 4'hF;
    S_A[62][1] = 4'hF;
    S_A[63][1] = 4'hF;
    S_A[64][1] = 4'hF;
    S_A[65][1] = 4'hF;
    S_A[66][1] = 4'hF;
    S_A[67][1] = 4'hF;
    S_A[68][1] = 4'hF;
    S_A[69][1] = 4'hF;
    S_A[70][1] = 4'hF;
    S_A[71][1] = 4'hF;
    S_A[72][1] = 4'hF;
    S_A[73][1] = 4'hF;
    S_A[74][1] = 4'hF;
    S_A[75][1] = 4'hF;
    S_A[76][1] = 4'hF;
    S_A[77][1] = 4'hF;
    S_A[78][1] = 4'hF;
    S_A[79][1] = 4'hF;
    S_A[80][1] = 4'hF;
    S_A[81][1] = 4'hF;
    S_A[82][1] = 4'hF;
    S_A[83][1] = 4'hF;
    S_A[84][1] = 4'hF;
    S_A[85][1] = 4'hF;
    S_A[86][1] = 4'hF;
    S_A[87][1] = 4'hF;
    S_A[88][1] = 4'hF;
    S_A[89][1] = 4'hF;
    S_A[90][1] = 4'hF;
    S_A[91][1] = 4'hF;
    S_A[92][1] = 4'hF;
    S_A[93][1] = 4'hF;
    S_A[94][1] = 4'hF;
    S_A[95][1] = 4'hF;
    S_A[96][1] = 4'hF;
    S_A[97][1] = 4'hF;
    S_A[98][1] = 4'hF;
    S_A[99][1] = 4'hF;
    S_A[100][1] = 4'hF;
    S_A[101][1] = 4'hF;
    S_A[102][1] = 4'hF;
    S_A[103][1] = 4'hF;
    S_A[104][1] = 4'hF;
    S_A[105][1] = 4'hF;
    S_A[106][1] = 4'hF;
    S_A[107][1] = 4'hF;
    S_A[108][1] = 4'hF;
    S_A[109][1] = 4'hF;
    S_A[110][1] = 4'hF;
    S_A[111][1] = 4'hF;
    S_A[112][1] = 4'hF;
    S_A[113][1] = 4'hF;
    S_A[114][1] = 4'hF;
    S_A[0][2] = 4'hF;
    S_A[1][2] = 4'hF;
    S_A[2][2] = 4'hF;
    S_A[3][2] = 4'hF;
    S_A[4][2] = 4'hF;
    S_A[5][2] = 4'hF;
    S_A[6][2] = 4'hF;
    S_A[7][2] = 4'hC;
    S_A[8][2] = 4'hC;
    S_A[9][2] = 4'hC;
    S_A[10][2] = 4'hC;
    S_A[11][2] = 4'hC;
    S_A[12][2] = 4'hC;
    S_A[13][2] = 4'hC;
    S_A[14][2] = 4'hC;
    S_A[15][2] = 4'hC;
    S_A[16][2] = 4'hC;
    S_A[17][2] = 4'hC;
    S_A[18][2] = 4'hC;
    S_A[19][2] = 4'hC;
    S_A[20][2] = 4'hC;
    S_A[21][2] = 4'hC;
    S_A[22][2] = 4'hF;
    S_A[23][2] = 4'hF;
    S_A[24][2] = 4'hF;
    S_A[25][2] = 4'hF;
    S_A[26][2] = 4'hF;
    S_A[27][2] = 4'hF;
    S_A[28][2] = 4'hF;
    S_A[29][2] = 4'hF;
    S_A[30][2] = 4'hF;
    S_A[31][2] = 4'hF;
    S_A[32][2] = 4'hF;
    S_A[33][2] = 4'hF;
    S_A[34][2] = 4'hF;
    S_A[35][2] = 4'hF;
    S_A[36][2] = 4'hF;
    S_A[37][2] = 4'hF;
    S_A[38][2] = 4'hF;
    S_A[39][2] = 4'hF;
    S_A[40][2] = 4'hF;
    S_A[41][2] = 4'hF;
    S_A[42][2] = 4'hF;
    S_A[43][2] = 4'hF;
    S_A[44][2] = 4'hF;
    S_A[45][2] = 4'hF;
    S_A[46][2] = 4'hF;
    S_A[47][2] = 4'hF;
    S_A[48][2] = 4'hF;
    S_A[49][2] = 4'hF;
    S_A[50][2] = 4'hF;
    S_A[51][2] = 4'hF;
    S_A[52][2] = 4'hF;
    S_A[53][2] = 4'hF;
    S_A[54][2] = 4'hF;
    S_A[55][2] = 4'hF;
    S_A[56][2] = 4'hF;
    S_A[57][2] = 4'hF;
    S_A[58][2] = 4'hF;
    S_A[59][2] = 4'hF;
    S_A[60][2] = 4'hF;
    S_A[61][2] = 4'hF;
    S_A[62][2] = 4'hF;
    S_A[63][2] = 4'hF;
    S_A[64][2] = 4'hF;
    S_A[65][2] = 4'hF;
    S_A[66][2] = 4'hF;
    S_A[67][2] = 4'hF;
    S_A[68][2] = 4'hF;
    S_A[69][2] = 4'hF;
    S_A[70][2] = 4'hF;
    S_A[71][2] = 4'hF;
    S_A[72][2] = 4'hF;
    S_A[73][2] = 4'hF;
    S_A[74][2] = 4'hF;
    S_A[75][2] = 4'hF;
    S_A[76][2] = 4'hF;
    S_A[77][2] = 4'hF;
    S_A[78][2] = 4'hF;
    S_A[79][2] = 4'hF;
    S_A[80][2] = 4'hF;
    S_A[81][2] = 4'hF;
    S_A[82][2] = 4'hF;
    S_A[83][2] = 4'hF;
    S_A[84][2] = 4'hF;
    S_A[85][2] = 4'hF;
    S_A[86][2] = 4'hF;
    S_A[87][2] = 4'hF;
    S_A[88][2] = 4'hF;
    S_A[89][2] = 4'hF;
    S_A[90][2] = 4'hF;
    S_A[91][2] = 4'hF;
    S_A[92][2] = 4'hF;
    S_A[93][2] = 4'hF;
    S_A[94][2] = 4'hF;
    S_A[95][2] = 4'hF;
    S_A[96][2] = 4'hF;
    S_A[97][2] = 4'hF;
    S_A[98][2] = 4'hF;
    S_A[99][2] = 4'hF;
    S_A[100][2] = 4'hF;
    S_A[101][2] = 4'hF;
    S_A[102][2] = 4'hF;
    S_A[103][2] = 4'hF;
    S_A[104][2] = 4'hF;
    S_A[105][2] = 4'hF;
    S_A[106][2] = 4'hF;
    S_A[107][2] = 4'hF;
    S_A[108][2] = 4'hF;
    S_A[109][2] = 4'hF;
    S_A[110][2] = 4'hF;
    S_A[111][2] = 4'hF;
    S_A[112][2] = 4'hF;
    S_A[113][2] = 4'hF;
    S_A[114][2] = 4'hF;
    S_A[0][3] = 4'hF;
    S_A[1][3] = 4'hF;
    S_A[2][3] = 4'hF;
    S_A[3][3] = 4'hF;
    S_A[4][3] = 4'hF;
    S_A[5][3] = 4'hF;
    S_A[6][3] = 4'hF;
    S_A[7][3] = 4'hC;
    S_A[8][3] = 4'hC;
    S_A[9][3] = 4'hC;
    S_A[10][3] = 4'hC;
    S_A[11][3] = 4'hC;
    S_A[12][3] = 4'hC;
    S_A[13][3] = 4'hC;
    S_A[14][3] = 4'hC;
    S_A[15][3] = 4'hC;
    S_A[16][3] = 4'hC;
    S_A[17][3] = 4'hC;
    S_A[18][3] = 4'hC;
    S_A[19][3] = 4'hC;
    S_A[20][3] = 4'hC;
    S_A[21][3] = 4'hC;
    S_A[22][3] = 4'hF;
    S_A[23][3] = 4'hF;
    S_A[24][3] = 4'hF;
    S_A[25][3] = 4'hF;
    S_A[26][3] = 4'hF;
    S_A[27][3] = 4'hF;
    S_A[28][3] = 4'hF;
    S_A[29][3] = 4'hF;
    S_A[30][3] = 4'hF;
    S_A[31][3] = 4'hF;
    S_A[32][3] = 4'hF;
    S_A[33][3] = 4'hF;
    S_A[34][3] = 4'hF;
    S_A[35][3] = 4'hF;
    S_A[36][3] = 4'hF;
    S_A[37][3] = 4'hF;
    S_A[38][3] = 4'hF;
    S_A[39][3] = 4'hF;
    S_A[40][3] = 4'hF;
    S_A[41][3] = 4'hF;
    S_A[42][3] = 4'hF;
    S_A[43][3] = 4'hF;
    S_A[44][3] = 4'hF;
    S_A[45][3] = 4'hF;
    S_A[46][3] = 4'hF;
    S_A[47][3] = 4'hF;
    S_A[48][3] = 4'hF;
    S_A[49][3] = 4'hF;
    S_A[50][3] = 4'hF;
    S_A[51][3] = 4'hF;
    S_A[52][3] = 4'hF;
    S_A[53][3] = 4'hF;
    S_A[54][3] = 4'hF;
    S_A[55][3] = 4'hF;
    S_A[56][3] = 4'hF;
    S_A[57][3] = 4'hF;
    S_A[58][3] = 4'hF;
    S_A[59][3] = 4'hF;
    S_A[60][3] = 4'hF;
    S_A[61][3] = 4'hF;
    S_A[62][3] = 4'hF;
    S_A[63][3] = 4'hF;
    S_A[64][3] = 4'hF;
    S_A[65][3] = 4'hF;
    S_A[66][3] = 4'hF;
    S_A[67][3] = 4'hF;
    S_A[68][3] = 4'hF;
    S_A[69][3] = 4'hF;
    S_A[70][3] = 4'hF;
    S_A[71][3] = 4'hF;
    S_A[72][3] = 4'hF;
    S_A[73][3] = 4'hF;
    S_A[74][3] = 4'hF;
    S_A[75][3] = 4'hF;
    S_A[76][3] = 4'hF;
    S_A[77][3] = 4'hF;
    S_A[78][3] = 4'hF;
    S_A[79][3] = 4'hF;
    S_A[80][3] = 4'hF;
    S_A[81][3] = 4'hF;
    S_A[82][3] = 4'hF;
    S_A[83][3] = 4'hF;
    S_A[84][3] = 4'hF;
    S_A[85][3] = 4'hF;
    S_A[86][3] = 4'hF;
    S_A[87][3] = 4'hF;
    S_A[88][3] = 4'hF;
    S_A[89][3] = 4'hF;
    S_A[90][3] = 4'hF;
    S_A[91][3] = 4'hF;
    S_A[92][3] = 4'hF;
    S_A[93][3] = 4'hF;
    S_A[94][3] = 4'hF;
    S_A[95][3] = 4'hF;
    S_A[96][3] = 4'hF;
    S_A[97][3] = 4'hF;
    S_A[98][3] = 4'hF;
    S_A[99][3] = 4'hF;
    S_A[100][3] = 4'hF;
    S_A[101][3] = 4'hF;
    S_A[102][3] = 4'hF;
    S_A[103][3] = 4'hF;
    S_A[104][3] = 4'hF;
    S_A[105][3] = 4'hF;
    S_A[106][3] = 4'hF;
    S_A[107][3] = 4'hF;
    S_A[108][3] = 4'hF;
    S_A[109][3] = 4'hF;
    S_A[110][3] = 4'hF;
    S_A[111][3] = 4'hF;
    S_A[112][3] = 4'hF;
    S_A[113][3] = 4'hF;
    S_A[114][3] = 4'hF;
    S_A[0][4] = 4'hF;
    S_A[1][4] = 4'hF;
    S_A[2][4] = 4'hF;
    S_A[3][4] = 4'hF;
    S_A[4][4] = 4'hF;
    S_A[5][4] = 4'hF;
    S_A[6][4] = 4'hF;
    S_A[7][4] = 4'hC;
    S_A[8][4] = 4'hC;
    S_A[9][4] = 4'hC;
    S_A[10][4] = 4'hC;
    S_A[11][4] = 4'hC;
    S_A[12][4] = 4'hC;
    S_A[13][4] = 4'hC;
    S_A[14][4] = 4'hC;
    S_A[15][4] = 4'hC;
    S_A[16][4] = 4'hC;
    S_A[17][4] = 4'hC;
    S_A[18][4] = 4'hC;
    S_A[19][4] = 4'hC;
    S_A[20][4] = 4'hC;
    S_A[21][4] = 4'hC;
    S_A[22][4] = 4'hF;
    S_A[23][4] = 4'hF;
    S_A[24][4] = 4'hF;
    S_A[25][4] = 4'hF;
    S_A[26][4] = 4'hF;
    S_A[27][4] = 4'hF;
    S_A[28][4] = 4'hF;
    S_A[29][4] = 4'hF;
    S_A[30][4] = 4'hF;
    S_A[31][4] = 4'hF;
    S_A[32][4] = 4'hF;
    S_A[33][4] = 4'hF;
    S_A[34][4] = 4'hF;
    S_A[35][4] = 4'hF;
    S_A[36][4] = 4'hF;
    S_A[37][4] = 4'hF;
    S_A[38][4] = 4'hF;
    S_A[39][4] = 4'hF;
    S_A[40][4] = 4'hF;
    S_A[41][4] = 4'hF;
    S_A[42][4] = 4'hF;
    S_A[43][4] = 4'hF;
    S_A[44][4] = 4'hF;
    S_A[45][4] = 4'hF;
    S_A[46][4] = 4'hF;
    S_A[47][4] = 4'hF;
    S_A[48][4] = 4'hF;
    S_A[49][4] = 4'hF;
    S_A[50][4] = 4'hF;
    S_A[51][4] = 4'hF;
    S_A[52][4] = 4'hF;
    S_A[53][4] = 4'hF;
    S_A[54][4] = 4'hF;
    S_A[55][4] = 4'hF;
    S_A[56][4] = 4'hF;
    S_A[57][4] = 4'hF;
    S_A[58][4] = 4'hF;
    S_A[59][4] = 4'hF;
    S_A[60][4] = 4'hF;
    S_A[61][4] = 4'hF;
    S_A[62][4] = 4'hF;
    S_A[63][4] = 4'hF;
    S_A[64][4] = 4'hF;
    S_A[65][4] = 4'hF;
    S_A[66][4] = 4'hF;
    S_A[67][4] = 4'hF;
    S_A[68][4] = 4'hF;
    S_A[69][4] = 4'hF;
    S_A[70][4] = 4'hF;
    S_A[71][4] = 4'hF;
    S_A[72][4] = 4'hF;
    S_A[73][4] = 4'hF;
    S_A[74][4] = 4'hF;
    S_A[75][4] = 4'hF;
    S_A[76][4] = 4'hF;
    S_A[77][4] = 4'hF;
    S_A[78][4] = 4'hF;
    S_A[79][4] = 4'hF;
    S_A[80][4] = 4'hF;
    S_A[81][4] = 4'hF;
    S_A[82][4] = 4'hF;
    S_A[83][4] = 4'hF;
    S_A[84][4] = 4'hF;
    S_A[85][4] = 4'hF;
    S_A[86][4] = 4'hF;
    S_A[87][4] = 4'hF;
    S_A[88][4] = 4'hF;
    S_A[89][4] = 4'hF;
    S_A[90][4] = 4'hF;
    S_A[91][4] = 4'hF;
    S_A[92][4] = 4'hF;
    S_A[93][4] = 4'hF;
    S_A[94][4] = 4'hF;
    S_A[95][4] = 4'hF;
    S_A[96][4] = 4'hF;
    S_A[97][4] = 4'hF;
    S_A[98][4] = 4'hF;
    S_A[99][4] = 4'hF;
    S_A[100][4] = 4'hF;
    S_A[101][4] = 4'hF;
    S_A[102][4] = 4'hF;
    S_A[103][4] = 4'hF;
    S_A[104][4] = 4'hF;
    S_A[105][4] = 4'hF;
    S_A[106][4] = 4'hF;
    S_A[107][4] = 4'hF;
    S_A[108][4] = 4'hF;
    S_A[109][4] = 4'hF;
    S_A[110][4] = 4'hF;
    S_A[111][4] = 4'hF;
    S_A[112][4] = 4'hF;
    S_A[113][4] = 4'hF;
    S_A[114][4] = 4'hF;
    S_A[0][5] = 4'hF;
    S_A[1][5] = 4'hF;
    S_A[2][5] = 4'hF;
    S_A[3][5] = 4'hF;
    S_A[4][5] = 4'hF;
    S_A[5][5] = 4'hF;
    S_A[6][5] = 4'hF;
    S_A[7][5] = 4'hC;
    S_A[8][5] = 4'hC;
    S_A[9][5] = 4'hC;
    S_A[10][5] = 4'hC;
    S_A[11][5] = 4'hC;
    S_A[12][5] = 4'hC;
    S_A[13][5] = 4'hC;
    S_A[14][5] = 4'hC;
    S_A[15][5] = 4'hC;
    S_A[16][5] = 4'hC;
    S_A[17][5] = 4'hC;
    S_A[18][5] = 4'hC;
    S_A[19][5] = 4'hC;
    S_A[20][5] = 4'hC;
    S_A[21][5] = 4'hC;
    S_A[22][5] = 4'hF;
    S_A[23][5] = 4'hF;
    S_A[24][5] = 4'hF;
    S_A[25][5] = 4'hF;
    S_A[26][5] = 4'hF;
    S_A[27][5] = 4'hF;
    S_A[28][5] = 4'hF;
    S_A[29][5] = 4'hF;
    S_A[30][5] = 4'hF;
    S_A[31][5] = 4'hF;
    S_A[32][5] = 4'hF;
    S_A[33][5] = 4'hF;
    S_A[34][5] = 4'hF;
    S_A[35][5] = 4'hF;
    S_A[36][5] = 4'hF;
    S_A[37][5] = 4'hF;
    S_A[38][5] = 4'hF;
    S_A[39][5] = 4'hF;
    S_A[40][5] = 4'hF;
    S_A[41][5] = 4'hF;
    S_A[42][5] = 4'hF;
    S_A[43][5] = 4'hF;
    S_A[44][5] = 4'hF;
    S_A[45][5] = 4'hF;
    S_A[46][5] = 4'hF;
    S_A[47][5] = 4'hF;
    S_A[48][5] = 4'hF;
    S_A[49][5] = 4'hF;
    S_A[50][5] = 4'hF;
    S_A[51][5] = 4'hF;
    S_A[52][5] = 4'hF;
    S_A[53][5] = 4'hF;
    S_A[54][5] = 4'hF;
    S_A[55][5] = 4'hF;
    S_A[56][5] = 4'hF;
    S_A[57][5] = 4'hF;
    S_A[58][5] = 4'hF;
    S_A[59][5] = 4'hF;
    S_A[60][5] = 4'hF;
    S_A[61][5] = 4'hF;
    S_A[62][5] = 4'hF;
    S_A[63][5] = 4'hF;
    S_A[64][5] = 4'hF;
    S_A[65][5] = 4'hF;
    S_A[66][5] = 4'hF;
    S_A[67][5] = 4'hF;
    S_A[68][5] = 4'hF;
    S_A[69][5] = 4'hF;
    S_A[70][5] = 4'hF;
    S_A[71][5] = 4'hF;
    S_A[72][5] = 4'hF;
    S_A[73][5] = 4'hF;
    S_A[74][5] = 4'hF;
    S_A[75][5] = 4'hF;
    S_A[76][5] = 4'hF;
    S_A[77][5] = 4'hF;
    S_A[78][5] = 4'hF;
    S_A[79][5] = 4'hF;
    S_A[80][5] = 4'hF;
    S_A[81][5] = 4'hF;
    S_A[82][5] = 4'hF;
    S_A[83][5] = 4'hF;
    S_A[84][5] = 4'hF;
    S_A[85][5] = 4'hF;
    S_A[86][5] = 4'hF;
    S_A[87][5] = 4'hF;
    S_A[88][5] = 4'hF;
    S_A[89][5] = 4'hF;
    S_A[90][5] = 4'hF;
    S_A[91][5] = 4'hF;
    S_A[92][5] = 4'hF;
    S_A[93][5] = 4'hF;
    S_A[94][5] = 4'hF;
    S_A[95][5] = 4'hF;
    S_A[96][5] = 4'hF;
    S_A[97][5] = 4'hF;
    S_A[98][5] = 4'hF;
    S_A[99][5] = 4'hF;
    S_A[100][5] = 4'hF;
    S_A[101][5] = 4'hF;
    S_A[102][5] = 4'hF;
    S_A[103][5] = 4'hF;
    S_A[104][5] = 4'hF;
    S_A[105][5] = 4'hF;
    S_A[106][5] = 4'hF;
    S_A[107][5] = 4'hF;
    S_A[108][5] = 4'hF;
    S_A[109][5] = 4'hF;
    S_A[110][5] = 4'hF;
    S_A[111][5] = 4'hF;
    S_A[112][5] = 4'hF;
    S_A[113][5] = 4'hF;
    S_A[114][5] = 4'hF;
    S_A[0][6] = 4'hF;
    S_A[1][6] = 4'hF;
    S_A[2][6] = 4'hF;
    S_A[3][6] = 4'hF;
    S_A[4][6] = 4'hF;
    S_A[5][6] = 4'hF;
    S_A[6][6] = 4'hF;
    S_A[7][6] = 4'hC;
    S_A[8][6] = 4'hC;
    S_A[9][6] = 4'hC;
    S_A[10][6] = 4'hC;
    S_A[11][6] = 4'hC;
    S_A[12][6] = 4'hC;
    S_A[13][6] = 4'hC;
    S_A[14][6] = 4'hC;
    S_A[15][6] = 4'hC;
    S_A[16][6] = 4'hC;
    S_A[17][6] = 4'hC;
    S_A[18][6] = 4'hC;
    S_A[19][6] = 4'hC;
    S_A[20][6] = 4'hC;
    S_A[21][6] = 4'hC;
    S_A[22][6] = 4'hF;
    S_A[23][6] = 4'hF;
    S_A[24][6] = 4'hF;
    S_A[25][6] = 4'hF;
    S_A[26][6] = 4'hF;
    S_A[27][6] = 4'hF;
    S_A[28][6] = 4'hF;
    S_A[29][6] = 4'hF;
    S_A[30][6] = 4'hF;
    S_A[31][6] = 4'hF;
    S_A[32][6] = 4'hF;
    S_A[33][6] = 4'hF;
    S_A[34][6] = 4'hF;
    S_A[35][6] = 4'hF;
    S_A[36][6] = 4'hF;
    S_A[37][6] = 4'hF;
    S_A[38][6] = 4'hF;
    S_A[39][6] = 4'hF;
    S_A[40][6] = 4'hF;
    S_A[41][6] = 4'hF;
    S_A[42][6] = 4'hF;
    S_A[43][6] = 4'hF;
    S_A[44][6] = 4'hF;
    S_A[45][6] = 4'hF;
    S_A[46][6] = 4'hF;
    S_A[47][6] = 4'hF;
    S_A[48][6] = 4'hF;
    S_A[49][6] = 4'hF;
    S_A[50][6] = 4'hF;
    S_A[51][6] = 4'hF;
    S_A[52][6] = 4'hF;
    S_A[53][6] = 4'hF;
    S_A[54][6] = 4'hF;
    S_A[55][6] = 4'hF;
    S_A[56][6] = 4'hF;
    S_A[57][6] = 4'hF;
    S_A[58][6] = 4'hF;
    S_A[59][6] = 4'hF;
    S_A[60][6] = 4'hF;
    S_A[61][6] = 4'hF;
    S_A[62][6] = 4'hF;
    S_A[63][6] = 4'hF;
    S_A[64][6] = 4'hF;
    S_A[65][6] = 4'hF;
    S_A[66][6] = 4'hF;
    S_A[67][6] = 4'hF;
    S_A[68][6] = 4'hF;
    S_A[69][6] = 4'hF;
    S_A[70][6] = 4'hF;
    S_A[71][6] = 4'hF;
    S_A[72][6] = 4'hF;
    S_A[73][6] = 4'hF;
    S_A[74][6] = 4'hF;
    S_A[75][6] = 4'hF;
    S_A[76][6] = 4'hF;
    S_A[77][6] = 4'hF;
    S_A[78][6] = 4'hF;
    S_A[79][6] = 4'hF;
    S_A[80][6] = 4'hF;
    S_A[81][6] = 4'hF;
    S_A[82][6] = 4'hF;
    S_A[83][6] = 4'hF;
    S_A[84][6] = 4'hF;
    S_A[85][6] = 4'hF;
    S_A[86][6] = 4'hF;
    S_A[87][6] = 4'hF;
    S_A[88][6] = 4'hF;
    S_A[89][6] = 4'hF;
    S_A[90][6] = 4'hF;
    S_A[91][6] = 4'hF;
    S_A[92][6] = 4'hF;
    S_A[93][6] = 4'hF;
    S_A[94][6] = 4'hF;
    S_A[95][6] = 4'hF;
    S_A[96][6] = 4'hF;
    S_A[97][6] = 4'hF;
    S_A[98][6] = 4'hF;
    S_A[99][6] = 4'hF;
    S_A[100][6] = 4'hF;
    S_A[101][6] = 4'hF;
    S_A[102][6] = 4'hF;
    S_A[103][6] = 4'hF;
    S_A[104][6] = 4'hF;
    S_A[105][6] = 4'hF;
    S_A[106][6] = 4'hF;
    S_A[107][6] = 4'hF;
    S_A[108][6] = 4'hF;
    S_A[109][6] = 4'hF;
    S_A[110][6] = 4'hF;
    S_A[111][6] = 4'hF;
    S_A[112][6] = 4'hF;
    S_A[113][6] = 4'hF;
    S_A[114][6] = 4'hF;
    S_A[0][7] = 4'hF;
    S_A[1][7] = 4'hF;
    S_A[2][7] = 4'hC;
    S_A[3][7] = 4'hC;
    S_A[4][7] = 4'hC;
    S_A[5][7] = 4'hC;
    S_A[6][7] = 4'hC;
    S_A[7][7] = 4'hF;
    S_A[8][7] = 4'hF;
    S_A[9][7] = 4'hF;
    S_A[10][7] = 4'hF;
    S_A[11][7] = 4'hF;
    S_A[12][7] = 4'hF;
    S_A[13][7] = 4'hF;
    S_A[14][7] = 4'hF;
    S_A[15][7] = 4'hF;
    S_A[16][7] = 4'hF;
    S_A[17][7] = 4'hF;
    S_A[18][7] = 4'hF;
    S_A[19][7] = 4'hF;
    S_A[20][7] = 4'hF;
    S_A[21][7] = 4'hF;
    S_A[22][7] = 4'hF;
    S_A[23][7] = 4'hF;
    S_A[24][7] = 4'hF;
    S_A[25][7] = 4'hF;
    S_A[26][7] = 4'hF;
    S_A[27][7] = 4'hF;
    S_A[28][7] = 4'hF;
    S_A[29][7] = 4'hF;
    S_A[30][7] = 4'hF;
    S_A[31][7] = 4'hF;
    S_A[32][7] = 4'hC;
    S_A[33][7] = 4'hC;
    S_A[34][7] = 4'hC;
    S_A[35][7] = 4'hC;
    S_A[36][7] = 4'hC;
    S_A[37][7] = 4'hC;
    S_A[38][7] = 4'hC;
    S_A[39][7] = 4'hC;
    S_A[40][7] = 4'hC;
    S_A[41][7] = 4'hC;
    S_A[42][7] = 4'hF;
    S_A[43][7] = 4'hF;
    S_A[44][7] = 4'hF;
    S_A[45][7] = 4'hF;
    S_A[46][7] = 4'hF;
    S_A[47][7] = 4'hF;
    S_A[48][7] = 4'hF;
    S_A[49][7] = 4'hF;
    S_A[50][7] = 4'hF;
    S_A[51][7] = 4'hF;
    S_A[52][7] = 4'hC;
    S_A[53][7] = 4'hC;
    S_A[54][7] = 4'hC;
    S_A[55][7] = 4'hC;
    S_A[56][7] = 4'hC;
    S_A[57][7] = 4'hC;
    S_A[58][7] = 4'hC;
    S_A[59][7] = 4'hC;
    S_A[60][7] = 4'hC;
    S_A[61][7] = 4'hC;
    S_A[62][7] = 4'hF;
    S_A[63][7] = 4'hF;
    S_A[64][7] = 4'hF;
    S_A[65][7] = 4'hF;
    S_A[66][7] = 4'hF;
    S_A[67][7] = 4'hF;
    S_A[68][7] = 4'hF;
    S_A[69][7] = 4'hF;
    S_A[70][7] = 4'hF;
    S_A[71][7] = 4'hF;
    S_A[72][7] = 4'hC;
    S_A[73][7] = 4'hC;
    S_A[74][7] = 4'hC;
    S_A[75][7] = 4'hC;
    S_A[76][7] = 4'hC;
    S_A[77][7] = 4'hF;
    S_A[78][7] = 4'hF;
    S_A[79][7] = 4'hF;
    S_A[80][7] = 4'hF;
    S_A[81][7] = 4'hF;
    S_A[82][7] = 4'hC;
    S_A[83][7] = 4'hC;
    S_A[84][7] = 4'hC;
    S_A[85][7] = 4'hC;
    S_A[86][7] = 4'hC;
    S_A[87][7] = 4'hF;
    S_A[88][7] = 4'hF;
    S_A[89][7] = 4'hF;
    S_A[90][7] = 4'hF;
    S_A[91][7] = 4'hF;
    S_A[92][7] = 4'hF;
    S_A[93][7] = 4'hF;
    S_A[94][7] = 4'hF;
    S_A[95][7] = 4'hF;
    S_A[96][7] = 4'hF;
    S_A[97][7] = 4'hC;
    S_A[98][7] = 4'hC;
    S_A[99][7] = 4'hC;
    S_A[100][7] = 4'hC;
    S_A[101][7] = 4'hC;
    S_A[102][7] = 4'hC;
    S_A[103][7] = 4'hC;
    S_A[104][7] = 4'hC;
    S_A[105][7] = 4'hC;
    S_A[106][7] = 4'hC;
    S_A[107][7] = 4'hF;
    S_A[108][7] = 4'hF;
    S_A[109][7] = 4'hF;
    S_A[110][7] = 4'hF;
    S_A[111][7] = 4'hF;
    S_A[112][7] = 4'hF;
    S_A[113][7] = 4'hF;
    S_A[114][7] = 4'hF;
    S_A[0][8] = 4'hF;
    S_A[1][8] = 4'hF;
    S_A[2][8] = 4'hC;
    S_A[3][8] = 4'hC;
    S_A[4][8] = 4'hC;
    S_A[5][8] = 4'hC;
    S_A[6][8] = 4'hC;
    S_A[7][8] = 4'hF;
    S_A[8][8] = 4'hF;
    S_A[9][8] = 4'hF;
    S_A[10][8] = 4'hF;
    S_A[11][8] = 4'hF;
    S_A[12][8] = 4'hF;
    S_A[13][8] = 4'hF;
    S_A[14][8] = 4'hF;
    S_A[15][8] = 4'hF;
    S_A[16][8] = 4'hF;
    S_A[17][8] = 4'hF;
    S_A[18][8] = 4'hF;
    S_A[19][8] = 4'hF;
    S_A[20][8] = 4'hF;
    S_A[21][8] = 4'hF;
    S_A[22][8] = 4'hF;
    S_A[23][8] = 4'hF;
    S_A[24][8] = 4'hF;
    S_A[25][8] = 4'hF;
    S_A[26][8] = 4'hF;
    S_A[27][8] = 4'hF;
    S_A[28][8] = 4'hF;
    S_A[29][8] = 4'hF;
    S_A[30][8] = 4'hF;
    S_A[31][8] = 4'hF;
    S_A[32][8] = 4'hC;
    S_A[33][8] = 4'hC;
    S_A[34][8] = 4'hC;
    S_A[35][8] = 4'hC;
    S_A[36][8] = 4'hC;
    S_A[37][8] = 4'hC;
    S_A[38][8] = 4'hC;
    S_A[39][8] = 4'hC;
    S_A[40][8] = 4'hC;
    S_A[41][8] = 4'hC;
    S_A[42][8] = 4'hF;
    S_A[43][8] = 4'hF;
    S_A[44][8] = 4'hF;
    S_A[45][8] = 4'hF;
    S_A[46][8] = 4'hF;
    S_A[47][8] = 4'hF;
    S_A[48][8] = 4'hF;
    S_A[49][8] = 4'hF;
    S_A[50][8] = 4'hF;
    S_A[51][8] = 4'hF;
    S_A[52][8] = 4'hC;
    S_A[53][8] = 4'hC;
    S_A[54][8] = 4'hC;
    S_A[55][8] = 4'hC;
    S_A[56][8] = 4'hC;
    S_A[57][8] = 4'hC;
    S_A[58][8] = 4'hC;
    S_A[59][8] = 4'hC;
    S_A[60][8] = 4'hC;
    S_A[61][8] = 4'hC;
    S_A[62][8] = 4'hF;
    S_A[63][8] = 4'hF;
    S_A[64][8] = 4'hF;
    S_A[65][8] = 4'hF;
    S_A[66][8] = 4'hF;
    S_A[67][8] = 4'hF;
    S_A[68][8] = 4'hF;
    S_A[69][8] = 4'hF;
    S_A[70][8] = 4'hF;
    S_A[71][8] = 4'hF;
    S_A[72][8] = 4'hC;
    S_A[73][8] = 4'hC;
    S_A[74][8] = 4'hC;
    S_A[75][8] = 4'hC;
    S_A[76][8] = 4'hC;
    S_A[77][8] = 4'hF;
    S_A[78][8] = 4'hF;
    S_A[79][8] = 4'hF;
    S_A[80][8] = 4'hF;
    S_A[81][8] = 4'hF;
    S_A[82][8] = 4'hC;
    S_A[83][8] = 4'hC;
    S_A[84][8] = 4'hC;
    S_A[85][8] = 4'hC;
    S_A[86][8] = 4'hC;
    S_A[87][8] = 4'hF;
    S_A[88][8] = 4'hF;
    S_A[89][8] = 4'hF;
    S_A[90][8] = 4'hF;
    S_A[91][8] = 4'hF;
    S_A[92][8] = 4'hF;
    S_A[93][8] = 4'hF;
    S_A[94][8] = 4'hF;
    S_A[95][8] = 4'hF;
    S_A[96][8] = 4'hF;
    S_A[97][8] = 4'hC;
    S_A[98][8] = 4'hC;
    S_A[99][8] = 4'hC;
    S_A[100][8] = 4'hC;
    S_A[101][8] = 4'hC;
    S_A[102][8] = 4'hC;
    S_A[103][8] = 4'hC;
    S_A[104][8] = 4'hC;
    S_A[105][8] = 4'hC;
    S_A[106][8] = 4'hC;
    S_A[107][8] = 4'hF;
    S_A[108][8] = 4'hF;
    S_A[109][8] = 4'hF;
    S_A[110][8] = 4'hF;
    S_A[111][8] = 4'hF;
    S_A[112][8] = 4'hF;
    S_A[113][8] = 4'hF;
    S_A[114][8] = 4'hF;
    S_A[0][9] = 4'hF;
    S_A[1][9] = 4'hF;
    S_A[2][9] = 4'hC;
    S_A[3][9] = 4'hC;
    S_A[4][9] = 4'hC;
    S_A[5][9] = 4'hC;
    S_A[6][9] = 4'hC;
    S_A[7][9] = 4'hF;
    S_A[8][9] = 4'hF;
    S_A[9][9] = 4'hF;
    S_A[10][9] = 4'hF;
    S_A[11][9] = 4'hF;
    S_A[12][9] = 4'hF;
    S_A[13][9] = 4'hF;
    S_A[14][9] = 4'hF;
    S_A[15][9] = 4'hF;
    S_A[16][9] = 4'hF;
    S_A[17][9] = 4'hF;
    S_A[18][9] = 4'hF;
    S_A[19][9] = 4'hF;
    S_A[20][9] = 4'hF;
    S_A[21][9] = 4'hF;
    S_A[22][9] = 4'hF;
    S_A[23][9] = 4'hF;
    S_A[24][9] = 4'hF;
    S_A[25][9] = 4'hF;
    S_A[26][9] = 4'hF;
    S_A[27][9] = 4'hF;
    S_A[28][9] = 4'hF;
    S_A[29][9] = 4'hF;
    S_A[30][9] = 4'hF;
    S_A[31][9] = 4'hF;
    S_A[32][9] = 4'hC;
    S_A[33][9] = 4'hC;
    S_A[34][9] = 4'hC;
    S_A[35][9] = 4'hC;
    S_A[36][9] = 4'hC;
    S_A[37][9] = 4'hC;
    S_A[38][9] = 4'hC;
    S_A[39][9] = 4'hC;
    S_A[40][9] = 4'hC;
    S_A[41][9] = 4'hC;
    S_A[42][9] = 4'hF;
    S_A[43][9] = 4'hF;
    S_A[44][9] = 4'hF;
    S_A[45][9] = 4'hF;
    S_A[46][9] = 4'hF;
    S_A[47][9] = 4'hF;
    S_A[48][9] = 4'hF;
    S_A[49][9] = 4'hF;
    S_A[50][9] = 4'hF;
    S_A[51][9] = 4'hF;
    S_A[52][9] = 4'hC;
    S_A[53][9] = 4'hC;
    S_A[54][9] = 4'hC;
    S_A[55][9] = 4'hC;
    S_A[56][9] = 4'hC;
    S_A[57][9] = 4'hC;
    S_A[58][9] = 4'hC;
    S_A[59][9] = 4'hC;
    S_A[60][9] = 4'hC;
    S_A[61][9] = 4'hC;
    S_A[62][9] = 4'hF;
    S_A[63][9] = 4'hF;
    S_A[64][9] = 4'hF;
    S_A[65][9] = 4'hF;
    S_A[66][9] = 4'hF;
    S_A[67][9] = 4'hF;
    S_A[68][9] = 4'hF;
    S_A[69][9] = 4'hF;
    S_A[70][9] = 4'hF;
    S_A[71][9] = 4'hF;
    S_A[72][9] = 4'hC;
    S_A[73][9] = 4'hC;
    S_A[74][9] = 4'hC;
    S_A[75][9] = 4'hC;
    S_A[76][9] = 4'hC;
    S_A[77][9] = 4'hF;
    S_A[78][9] = 4'hF;
    S_A[79][9] = 4'hF;
    S_A[80][9] = 4'hF;
    S_A[81][9] = 4'hF;
    S_A[82][9] = 4'hC;
    S_A[83][9] = 4'hC;
    S_A[84][9] = 4'hC;
    S_A[85][9] = 4'hC;
    S_A[86][9] = 4'hC;
    S_A[87][9] = 4'hF;
    S_A[88][9] = 4'hF;
    S_A[89][9] = 4'hF;
    S_A[90][9] = 4'hF;
    S_A[91][9] = 4'hF;
    S_A[92][9] = 4'hF;
    S_A[93][9] = 4'hF;
    S_A[94][9] = 4'hF;
    S_A[95][9] = 4'hF;
    S_A[96][9] = 4'hF;
    S_A[97][9] = 4'hC;
    S_A[98][9] = 4'hC;
    S_A[99][9] = 4'hC;
    S_A[100][9] = 4'hC;
    S_A[101][9] = 4'hC;
    S_A[102][9] = 4'hC;
    S_A[103][9] = 4'hC;
    S_A[104][9] = 4'hC;
    S_A[105][9] = 4'hC;
    S_A[106][9] = 4'hC;
    S_A[107][9] = 4'hF;
    S_A[108][9] = 4'hF;
    S_A[109][9] = 4'hF;
    S_A[110][9] = 4'hF;
    S_A[111][9] = 4'hF;
    S_A[112][9] = 4'hF;
    S_A[113][9] = 4'hF;
    S_A[114][9] = 4'hF;
    S_A[0][10] = 4'hF;
    S_A[1][10] = 4'hF;
    S_A[2][10] = 4'hC;
    S_A[3][10] = 4'hC;
    S_A[4][10] = 4'hC;
    S_A[5][10] = 4'hC;
    S_A[6][10] = 4'hC;
    S_A[7][10] = 4'hF;
    S_A[8][10] = 4'hF;
    S_A[9][10] = 4'hF;
    S_A[10][10] = 4'hF;
    S_A[11][10] = 4'hF;
    S_A[12][10] = 4'hF;
    S_A[13][10] = 4'hF;
    S_A[14][10] = 4'hF;
    S_A[15][10] = 4'hF;
    S_A[16][10] = 4'hF;
    S_A[17][10] = 4'hF;
    S_A[18][10] = 4'hF;
    S_A[19][10] = 4'hF;
    S_A[20][10] = 4'hF;
    S_A[21][10] = 4'hF;
    S_A[22][10] = 4'hF;
    S_A[23][10] = 4'hF;
    S_A[24][10] = 4'hF;
    S_A[25][10] = 4'hF;
    S_A[26][10] = 4'hF;
    S_A[27][10] = 4'hF;
    S_A[28][10] = 4'hF;
    S_A[29][10] = 4'hF;
    S_A[30][10] = 4'hF;
    S_A[31][10] = 4'hF;
    S_A[32][10] = 4'hC;
    S_A[33][10] = 4'hC;
    S_A[34][10] = 4'hC;
    S_A[35][10] = 4'hC;
    S_A[36][10] = 4'hC;
    S_A[37][10] = 4'hC;
    S_A[38][10] = 4'hC;
    S_A[39][10] = 4'hC;
    S_A[40][10] = 4'hC;
    S_A[41][10] = 4'hC;
    S_A[42][10] = 4'hF;
    S_A[43][10] = 4'hF;
    S_A[44][10] = 4'hF;
    S_A[45][10] = 4'hF;
    S_A[46][10] = 4'hF;
    S_A[47][10] = 4'hF;
    S_A[48][10] = 4'hF;
    S_A[49][10] = 4'hF;
    S_A[50][10] = 4'hF;
    S_A[51][10] = 4'hF;
    S_A[52][10] = 4'hC;
    S_A[53][10] = 4'hC;
    S_A[54][10] = 4'hC;
    S_A[55][10] = 4'hC;
    S_A[56][10] = 4'hC;
    S_A[57][10] = 4'hC;
    S_A[58][10] = 4'hC;
    S_A[59][10] = 4'hC;
    S_A[60][10] = 4'hC;
    S_A[61][10] = 4'hC;
    S_A[62][10] = 4'hF;
    S_A[63][10] = 4'hF;
    S_A[64][10] = 4'hF;
    S_A[65][10] = 4'hF;
    S_A[66][10] = 4'hF;
    S_A[67][10] = 4'hF;
    S_A[68][10] = 4'hF;
    S_A[69][10] = 4'hF;
    S_A[70][10] = 4'hF;
    S_A[71][10] = 4'hF;
    S_A[72][10] = 4'hC;
    S_A[73][10] = 4'hC;
    S_A[74][10] = 4'hC;
    S_A[75][10] = 4'hC;
    S_A[76][10] = 4'hC;
    S_A[77][10] = 4'hF;
    S_A[78][10] = 4'hF;
    S_A[79][10] = 4'hF;
    S_A[80][10] = 4'hF;
    S_A[81][10] = 4'hF;
    S_A[82][10] = 4'hC;
    S_A[83][10] = 4'hC;
    S_A[84][10] = 4'hC;
    S_A[85][10] = 4'hC;
    S_A[86][10] = 4'hC;
    S_A[87][10] = 4'hF;
    S_A[88][10] = 4'hF;
    S_A[89][10] = 4'hF;
    S_A[90][10] = 4'hF;
    S_A[91][10] = 4'hF;
    S_A[92][10] = 4'hF;
    S_A[93][10] = 4'hF;
    S_A[94][10] = 4'hF;
    S_A[95][10] = 4'hF;
    S_A[96][10] = 4'hF;
    S_A[97][10] = 4'hC;
    S_A[98][10] = 4'hC;
    S_A[99][10] = 4'hC;
    S_A[100][10] = 4'hC;
    S_A[101][10] = 4'hC;
    S_A[102][10] = 4'hC;
    S_A[103][10] = 4'hC;
    S_A[104][10] = 4'hC;
    S_A[105][10] = 4'hC;
    S_A[106][10] = 4'hC;
    S_A[107][10] = 4'hF;
    S_A[108][10] = 4'hF;
    S_A[109][10] = 4'hF;
    S_A[110][10] = 4'hF;
    S_A[111][10] = 4'hF;
    S_A[112][10] = 4'hF;
    S_A[113][10] = 4'hF;
    S_A[114][10] = 4'hF;
    S_A[0][11] = 4'hF;
    S_A[1][11] = 4'hF;
    S_A[2][11] = 4'hC;
    S_A[3][11] = 4'hC;
    S_A[4][11] = 4'hC;
    S_A[5][11] = 4'hC;
    S_A[6][11] = 4'hC;
    S_A[7][11] = 4'hF;
    S_A[8][11] = 4'hF;
    S_A[9][11] = 4'hF;
    S_A[10][11] = 4'hF;
    S_A[11][11] = 4'hF;
    S_A[12][11] = 4'hF;
    S_A[13][11] = 4'hF;
    S_A[14][11] = 4'hF;
    S_A[15][11] = 4'hF;
    S_A[16][11] = 4'hF;
    S_A[17][11] = 4'hF;
    S_A[18][11] = 4'hF;
    S_A[19][11] = 4'hF;
    S_A[20][11] = 4'hF;
    S_A[21][11] = 4'hF;
    S_A[22][11] = 4'hF;
    S_A[23][11] = 4'hF;
    S_A[24][11] = 4'hF;
    S_A[25][11] = 4'hF;
    S_A[26][11] = 4'hF;
    S_A[27][11] = 4'hF;
    S_A[28][11] = 4'hF;
    S_A[29][11] = 4'hF;
    S_A[30][11] = 4'hF;
    S_A[31][11] = 4'hF;
    S_A[32][11] = 4'hC;
    S_A[33][11] = 4'hC;
    S_A[34][11] = 4'hC;
    S_A[35][11] = 4'hC;
    S_A[36][11] = 4'hC;
    S_A[37][11] = 4'hC;
    S_A[38][11] = 4'hC;
    S_A[39][11] = 4'hC;
    S_A[40][11] = 4'hC;
    S_A[41][11] = 4'hC;
    S_A[42][11] = 4'hF;
    S_A[43][11] = 4'hF;
    S_A[44][11] = 4'hF;
    S_A[45][11] = 4'hF;
    S_A[46][11] = 4'hF;
    S_A[47][11] = 4'hF;
    S_A[48][11] = 4'hF;
    S_A[49][11] = 4'hF;
    S_A[50][11] = 4'hF;
    S_A[51][11] = 4'hF;
    S_A[52][11] = 4'hC;
    S_A[53][11] = 4'hC;
    S_A[54][11] = 4'hC;
    S_A[55][11] = 4'hC;
    S_A[56][11] = 4'hC;
    S_A[57][11] = 4'hC;
    S_A[58][11] = 4'hC;
    S_A[59][11] = 4'hC;
    S_A[60][11] = 4'hC;
    S_A[61][11] = 4'hC;
    S_A[62][11] = 4'hF;
    S_A[63][11] = 4'hF;
    S_A[64][11] = 4'hF;
    S_A[65][11] = 4'hF;
    S_A[66][11] = 4'hF;
    S_A[67][11] = 4'hF;
    S_A[68][11] = 4'hF;
    S_A[69][11] = 4'hF;
    S_A[70][11] = 4'hF;
    S_A[71][11] = 4'hF;
    S_A[72][11] = 4'hC;
    S_A[73][11] = 4'hC;
    S_A[74][11] = 4'hC;
    S_A[75][11] = 4'hC;
    S_A[76][11] = 4'hC;
    S_A[77][11] = 4'hF;
    S_A[78][11] = 4'hF;
    S_A[79][11] = 4'hF;
    S_A[80][11] = 4'hF;
    S_A[81][11] = 4'hF;
    S_A[82][11] = 4'hC;
    S_A[83][11] = 4'hC;
    S_A[84][11] = 4'hC;
    S_A[85][11] = 4'hC;
    S_A[86][11] = 4'hC;
    S_A[87][11] = 4'hF;
    S_A[88][11] = 4'hF;
    S_A[89][11] = 4'hF;
    S_A[90][11] = 4'hF;
    S_A[91][11] = 4'hF;
    S_A[92][11] = 4'hF;
    S_A[93][11] = 4'hF;
    S_A[94][11] = 4'hF;
    S_A[95][11] = 4'hF;
    S_A[96][11] = 4'hF;
    S_A[97][11] = 4'hC;
    S_A[98][11] = 4'hC;
    S_A[99][11] = 4'hC;
    S_A[100][11] = 4'hC;
    S_A[101][11] = 4'hC;
    S_A[102][11] = 4'hC;
    S_A[103][11] = 4'hC;
    S_A[104][11] = 4'hC;
    S_A[105][11] = 4'hC;
    S_A[106][11] = 4'hC;
    S_A[107][11] = 4'hF;
    S_A[108][11] = 4'hF;
    S_A[109][11] = 4'hF;
    S_A[110][11] = 4'hF;
    S_A[111][11] = 4'hF;
    S_A[112][11] = 4'hF;
    S_A[113][11] = 4'hF;
    S_A[114][11] = 4'hF;
    S_A[0][12] = 4'hF;
    S_A[1][12] = 4'hF;
    S_A[2][12] = 4'hF;
    S_A[3][12] = 4'hF;
    S_A[4][12] = 4'hF;
    S_A[5][12] = 4'hF;
    S_A[6][12] = 4'hF;
    S_A[7][12] = 4'hC;
    S_A[8][12] = 4'hC;
    S_A[9][12] = 4'hC;
    S_A[10][12] = 4'hC;
    S_A[11][12] = 4'hC;
    S_A[12][12] = 4'hC;
    S_A[13][12] = 4'hC;
    S_A[14][12] = 4'hC;
    S_A[15][12] = 4'hC;
    S_A[16][12] = 4'hC;
    S_A[17][12] = 4'hF;
    S_A[18][12] = 4'hF;
    S_A[19][12] = 4'hF;
    S_A[20][12] = 4'hF;
    S_A[21][12] = 4'hF;
    S_A[22][12] = 4'hF;
    S_A[23][12] = 4'hF;
    S_A[24][12] = 4'hF;
    S_A[25][12] = 4'hF;
    S_A[26][12] = 4'hF;
    S_A[27][12] = 4'hC;
    S_A[28][12] = 4'hC;
    S_A[29][12] = 4'hC;
    S_A[30][12] = 4'hC;
    S_A[31][12] = 4'hC;
    S_A[32][12] = 4'hF;
    S_A[33][12] = 4'hF;
    S_A[34][12] = 4'hF;
    S_A[35][12] = 4'hF;
    S_A[36][12] = 4'hF;
    S_A[37][12] = 4'hF;
    S_A[38][12] = 4'hF;
    S_A[39][12] = 4'hF;
    S_A[40][12] = 4'hF;
    S_A[41][12] = 4'hF;
    S_A[42][12] = 4'hF;
    S_A[43][12] = 4'hF;
    S_A[44][12] = 4'hF;
    S_A[45][12] = 4'hF;
    S_A[46][12] = 4'hF;
    S_A[47][12] = 4'hC;
    S_A[48][12] = 4'hC;
    S_A[49][12] = 4'hC;
    S_A[50][12] = 4'hC;
    S_A[51][12] = 4'hC;
    S_A[52][12] = 4'hF;
    S_A[53][12] = 4'hF;
    S_A[54][12] = 4'hF;
    S_A[55][12] = 4'hF;
    S_A[56][12] = 4'hF;
    S_A[57][12] = 4'hF;
    S_A[58][12] = 4'hF;
    S_A[59][12] = 4'hF;
    S_A[60][12] = 4'hF;
    S_A[61][12] = 4'hF;
    S_A[62][12] = 4'hC;
    S_A[63][12] = 4'hC;
    S_A[64][12] = 4'hC;
    S_A[65][12] = 4'hC;
    S_A[66][12] = 4'hC;
    S_A[67][12] = 4'hF;
    S_A[68][12] = 4'hF;
    S_A[69][12] = 4'hF;
    S_A[70][12] = 4'hF;
    S_A[71][12] = 4'hF;
    S_A[72][12] = 4'hC;
    S_A[73][12] = 4'hC;
    S_A[74][12] = 4'hC;
    S_A[75][12] = 4'hC;
    S_A[76][12] = 4'hC;
    S_A[77][12] = 4'hC;
    S_A[78][12] = 4'hC;
    S_A[79][12] = 4'hC;
    S_A[80][12] = 4'hC;
    S_A[81][12] = 4'hC;
    S_A[82][12] = 4'hF;
    S_A[83][12] = 4'hF;
    S_A[84][12] = 4'hF;
    S_A[85][12] = 4'hF;
    S_A[86][12] = 4'hF;
    S_A[87][12] = 4'hF;
    S_A[88][12] = 4'hF;
    S_A[89][12] = 4'hF;
    S_A[90][12] = 4'hF;
    S_A[91][12] = 4'hF;
    S_A[92][12] = 4'hC;
    S_A[93][12] = 4'hC;
    S_A[94][12] = 4'hC;
    S_A[95][12] = 4'hC;
    S_A[96][12] = 4'hC;
    S_A[97][12] = 4'hF;
    S_A[98][12] = 4'hF;
    S_A[99][12] = 4'hF;
    S_A[100][12] = 4'hF;
    S_A[101][12] = 4'hF;
    S_A[102][12] = 4'hC;
    S_A[103][12] = 4'hC;
    S_A[104][12] = 4'hC;
    S_A[105][12] = 4'hC;
    S_A[106][12] = 4'hC;
    S_A[107][12] = 4'hC;
    S_A[108][12] = 4'hC;
    S_A[109][12] = 4'hC;
    S_A[110][12] = 4'hC;
    S_A[111][12] = 4'hC;
    S_A[112][12] = 4'hF;
    S_A[113][12] = 4'hF;
    S_A[114][12] = 4'hF;
    S_A[0][13] = 4'hF;
    S_A[1][13] = 4'hF;
    S_A[2][13] = 4'hF;
    S_A[3][13] = 4'hF;
    S_A[4][13] = 4'hF;
    S_A[5][13] = 4'hF;
    S_A[6][13] = 4'hF;
    S_A[7][13] = 4'hC;
    S_A[8][13] = 4'hC;
    S_A[9][13] = 4'hC;
    S_A[10][13] = 4'hC;
    S_A[11][13] = 4'hC;
    S_A[12][13] = 4'hC;
    S_A[13][13] = 4'hC;
    S_A[14][13] = 4'hC;
    S_A[15][13] = 4'hC;
    S_A[16][13] = 4'hC;
    S_A[17][13] = 4'hF;
    S_A[18][13] = 4'hF;
    S_A[19][13] = 4'hF;
    S_A[20][13] = 4'hF;
    S_A[21][13] = 4'hF;
    S_A[22][13] = 4'hF;
    S_A[23][13] = 4'hF;
    S_A[24][13] = 4'hF;
    S_A[25][13] = 4'hF;
    S_A[26][13] = 4'hF;
    S_A[27][13] = 4'hC;
    S_A[28][13] = 4'hC;
    S_A[29][13] = 4'hC;
    S_A[30][13] = 4'hC;
    S_A[31][13] = 4'hC;
    S_A[32][13] = 4'hF;
    S_A[33][13] = 4'hF;
    S_A[34][13] = 4'hF;
    S_A[35][13] = 4'hF;
    S_A[36][13] = 4'hF;
    S_A[37][13] = 4'hF;
    S_A[38][13] = 4'hF;
    S_A[39][13] = 4'hF;
    S_A[40][13] = 4'hF;
    S_A[41][13] = 4'hF;
    S_A[42][13] = 4'hF;
    S_A[43][13] = 4'hF;
    S_A[44][13] = 4'hF;
    S_A[45][13] = 4'hF;
    S_A[46][13] = 4'hF;
    S_A[47][13] = 4'hC;
    S_A[48][13] = 4'hC;
    S_A[49][13] = 4'hC;
    S_A[50][13] = 4'hC;
    S_A[51][13] = 4'hC;
    S_A[52][13] = 4'hF;
    S_A[53][13] = 4'hF;
    S_A[54][13] = 4'hF;
    S_A[55][13] = 4'hF;
    S_A[56][13] = 4'hF;
    S_A[57][13] = 4'hF;
    S_A[58][13] = 4'hF;
    S_A[59][13] = 4'hF;
    S_A[60][13] = 4'hF;
    S_A[61][13] = 4'hF;
    S_A[62][13] = 4'hC;
    S_A[63][13] = 4'hC;
    S_A[64][13] = 4'hC;
    S_A[65][13] = 4'hC;
    S_A[66][13] = 4'hC;
    S_A[67][13] = 4'hF;
    S_A[68][13] = 4'hF;
    S_A[69][13] = 4'hF;
    S_A[70][13] = 4'hF;
    S_A[71][13] = 4'hF;
    S_A[72][13] = 4'hC;
    S_A[73][13] = 4'hC;
    S_A[74][13] = 4'hC;
    S_A[75][13] = 4'hC;
    S_A[76][13] = 4'hC;
    S_A[77][13] = 4'hC;
    S_A[78][13] = 4'hC;
    S_A[79][13] = 4'hC;
    S_A[80][13] = 4'hC;
    S_A[81][13] = 4'hC;
    S_A[82][13] = 4'hF;
    S_A[83][13] = 4'hF;
    S_A[84][13] = 4'hF;
    S_A[85][13] = 4'hF;
    S_A[86][13] = 4'hF;
    S_A[87][13] = 4'hF;
    S_A[88][13] = 4'hF;
    S_A[89][13] = 4'hF;
    S_A[90][13] = 4'hF;
    S_A[91][13] = 4'hF;
    S_A[92][13] = 4'hC;
    S_A[93][13] = 4'hC;
    S_A[94][13] = 4'hC;
    S_A[95][13] = 4'hC;
    S_A[96][13] = 4'hC;
    S_A[97][13] = 4'hF;
    S_A[98][13] = 4'hF;
    S_A[99][13] = 4'hF;
    S_A[100][13] = 4'hF;
    S_A[101][13] = 4'hF;
    S_A[102][13] = 4'hC;
    S_A[103][13] = 4'hC;
    S_A[104][13] = 4'hC;
    S_A[105][13] = 4'hC;
    S_A[106][13] = 4'hC;
    S_A[107][13] = 4'hC;
    S_A[108][13] = 4'hC;
    S_A[109][13] = 4'hC;
    S_A[110][13] = 4'hC;
    S_A[111][13] = 4'hC;
    S_A[112][13] = 4'hF;
    S_A[113][13] = 4'hF;
    S_A[114][13] = 4'hF;
    S_A[0][14] = 4'hF;
    S_A[1][14] = 4'hF;
    S_A[2][14] = 4'hF;
    S_A[3][14] = 4'hF;
    S_A[4][14] = 4'hF;
    S_A[5][14] = 4'hF;
    S_A[6][14] = 4'hF;
    S_A[7][14] = 4'hC;
    S_A[8][14] = 4'hC;
    S_A[9][14] = 4'hC;
    S_A[10][14] = 4'hC;
    S_A[11][14] = 4'hC;
    S_A[12][14] = 4'hC;
    S_A[13][14] = 4'hC;
    S_A[14][14] = 4'hC;
    S_A[15][14] = 4'hC;
    S_A[16][14] = 4'hC;
    S_A[17][14] = 4'hF;
    S_A[18][14] = 4'hF;
    S_A[19][14] = 4'hF;
    S_A[20][14] = 4'hF;
    S_A[21][14] = 4'hF;
    S_A[22][14] = 4'hF;
    S_A[23][14] = 4'hF;
    S_A[24][14] = 4'hF;
    S_A[25][14] = 4'hF;
    S_A[26][14] = 4'hF;
    S_A[27][14] = 4'hC;
    S_A[28][14] = 4'hC;
    S_A[29][14] = 4'hC;
    S_A[30][14] = 4'hC;
    S_A[31][14] = 4'hC;
    S_A[32][14] = 4'hF;
    S_A[33][14] = 4'hF;
    S_A[34][14] = 4'hF;
    S_A[35][14] = 4'hF;
    S_A[36][14] = 4'hF;
    S_A[37][14] = 4'hF;
    S_A[38][14] = 4'hF;
    S_A[39][14] = 4'hF;
    S_A[40][14] = 4'hF;
    S_A[41][14] = 4'hF;
    S_A[42][14] = 4'hF;
    S_A[43][14] = 4'hF;
    S_A[44][14] = 4'hF;
    S_A[45][14] = 4'hF;
    S_A[46][14] = 4'hF;
    S_A[47][14] = 4'hC;
    S_A[48][14] = 4'hC;
    S_A[49][14] = 4'hC;
    S_A[50][14] = 4'hC;
    S_A[51][14] = 4'hC;
    S_A[52][14] = 4'hF;
    S_A[53][14] = 4'hF;
    S_A[54][14] = 4'hF;
    S_A[55][14] = 4'hF;
    S_A[56][14] = 4'hF;
    S_A[57][14] = 4'hF;
    S_A[58][14] = 4'hF;
    S_A[59][14] = 4'hF;
    S_A[60][14] = 4'hF;
    S_A[61][14] = 4'hF;
    S_A[62][14] = 4'hC;
    S_A[63][14] = 4'hC;
    S_A[64][14] = 4'hC;
    S_A[65][14] = 4'hC;
    S_A[66][14] = 4'hC;
    S_A[67][14] = 4'hF;
    S_A[68][14] = 4'hF;
    S_A[69][14] = 4'hF;
    S_A[70][14] = 4'hF;
    S_A[71][14] = 4'hF;
    S_A[72][14] = 4'hC;
    S_A[73][14] = 4'hC;
    S_A[74][14] = 4'hC;
    S_A[75][14] = 4'hC;
    S_A[76][14] = 4'hC;
    S_A[77][14] = 4'hC;
    S_A[78][14] = 4'hC;
    S_A[79][14] = 4'hC;
    S_A[80][14] = 4'hC;
    S_A[81][14] = 4'hC;
    S_A[82][14] = 4'hF;
    S_A[83][14] = 4'hF;
    S_A[84][14] = 4'hF;
    S_A[85][14] = 4'hF;
    S_A[86][14] = 4'hF;
    S_A[87][14] = 4'hF;
    S_A[88][14] = 4'hF;
    S_A[89][14] = 4'hF;
    S_A[90][14] = 4'hF;
    S_A[91][14] = 4'hF;
    S_A[92][14] = 4'hC;
    S_A[93][14] = 4'hC;
    S_A[94][14] = 4'hC;
    S_A[95][14] = 4'hC;
    S_A[96][14] = 4'hC;
    S_A[97][14] = 4'hF;
    S_A[98][14] = 4'hF;
    S_A[99][14] = 4'hF;
    S_A[100][14] = 4'hF;
    S_A[101][14] = 4'hF;
    S_A[102][14] = 4'hC;
    S_A[103][14] = 4'hC;
    S_A[104][14] = 4'hC;
    S_A[105][14] = 4'hC;
    S_A[106][14] = 4'hC;
    S_A[107][14] = 4'hC;
    S_A[108][14] = 4'hC;
    S_A[109][14] = 4'hC;
    S_A[110][14] = 4'hC;
    S_A[111][14] = 4'hC;
    S_A[112][14] = 4'hF;
    S_A[113][14] = 4'hF;
    S_A[114][14] = 4'hF;
    S_A[0][15] = 4'hF;
    S_A[1][15] = 4'hF;
    S_A[2][15] = 4'hF;
    S_A[3][15] = 4'hF;
    S_A[4][15] = 4'hF;
    S_A[5][15] = 4'hF;
    S_A[6][15] = 4'hF;
    S_A[7][15] = 4'hC;
    S_A[8][15] = 4'hC;
    S_A[9][15] = 4'hC;
    S_A[10][15] = 4'hC;
    S_A[11][15] = 4'hC;
    S_A[12][15] = 4'hC;
    S_A[13][15] = 4'hC;
    S_A[14][15] = 4'hC;
    S_A[15][15] = 4'hC;
    S_A[16][15] = 4'hC;
    S_A[17][15] = 4'hF;
    S_A[18][15] = 4'hF;
    S_A[19][15] = 4'hF;
    S_A[20][15] = 4'hF;
    S_A[21][15] = 4'hF;
    S_A[22][15] = 4'hF;
    S_A[23][15] = 4'hF;
    S_A[24][15] = 4'hF;
    S_A[25][15] = 4'hF;
    S_A[26][15] = 4'hF;
    S_A[27][15] = 4'hC;
    S_A[28][15] = 4'hC;
    S_A[29][15] = 4'hC;
    S_A[30][15] = 4'hC;
    S_A[31][15] = 4'hC;
    S_A[32][15] = 4'hF;
    S_A[33][15] = 4'hF;
    S_A[34][15] = 4'hF;
    S_A[35][15] = 4'hF;
    S_A[36][15] = 4'hF;
    S_A[37][15] = 4'hF;
    S_A[38][15] = 4'hF;
    S_A[39][15] = 4'hF;
    S_A[40][15] = 4'hF;
    S_A[41][15] = 4'hF;
    S_A[42][15] = 4'hF;
    S_A[43][15] = 4'hF;
    S_A[44][15] = 4'hF;
    S_A[45][15] = 4'hF;
    S_A[46][15] = 4'hF;
    S_A[47][15] = 4'hC;
    S_A[48][15] = 4'hC;
    S_A[49][15] = 4'hC;
    S_A[50][15] = 4'hC;
    S_A[51][15] = 4'hC;
    S_A[52][15] = 4'hF;
    S_A[53][15] = 4'hF;
    S_A[54][15] = 4'hF;
    S_A[55][15] = 4'hF;
    S_A[56][15] = 4'hF;
    S_A[57][15] = 4'hF;
    S_A[58][15] = 4'hF;
    S_A[59][15] = 4'hF;
    S_A[60][15] = 4'hF;
    S_A[61][15] = 4'hF;
    S_A[62][15] = 4'hC;
    S_A[63][15] = 4'hC;
    S_A[64][15] = 4'hC;
    S_A[65][15] = 4'hC;
    S_A[66][15] = 4'hC;
    S_A[67][15] = 4'hF;
    S_A[68][15] = 4'hF;
    S_A[69][15] = 4'hF;
    S_A[70][15] = 4'hF;
    S_A[71][15] = 4'hF;
    S_A[72][15] = 4'hC;
    S_A[73][15] = 4'hC;
    S_A[74][15] = 4'hC;
    S_A[75][15] = 4'hC;
    S_A[76][15] = 4'hC;
    S_A[77][15] = 4'hC;
    S_A[78][15] = 4'hC;
    S_A[79][15] = 4'hC;
    S_A[80][15] = 4'hC;
    S_A[81][15] = 4'hC;
    S_A[82][15] = 4'hF;
    S_A[83][15] = 4'hF;
    S_A[84][15] = 4'hF;
    S_A[85][15] = 4'hF;
    S_A[86][15] = 4'hF;
    S_A[87][15] = 4'hF;
    S_A[88][15] = 4'hF;
    S_A[89][15] = 4'hF;
    S_A[90][15] = 4'hF;
    S_A[91][15] = 4'hF;
    S_A[92][15] = 4'hC;
    S_A[93][15] = 4'hC;
    S_A[94][15] = 4'hC;
    S_A[95][15] = 4'hC;
    S_A[96][15] = 4'hC;
    S_A[97][15] = 4'hF;
    S_A[98][15] = 4'hF;
    S_A[99][15] = 4'hF;
    S_A[100][15] = 4'hF;
    S_A[101][15] = 4'hF;
    S_A[102][15] = 4'hC;
    S_A[103][15] = 4'hC;
    S_A[104][15] = 4'hC;
    S_A[105][15] = 4'hC;
    S_A[106][15] = 4'hC;
    S_A[107][15] = 4'hC;
    S_A[108][15] = 4'hC;
    S_A[109][15] = 4'hC;
    S_A[110][15] = 4'hC;
    S_A[111][15] = 4'hC;
    S_A[112][15] = 4'hF;
    S_A[113][15] = 4'hF;
    S_A[114][15] = 4'hF;
    S_A[0][16] = 4'hF;
    S_A[1][16] = 4'hF;
    S_A[2][16] = 4'hF;
    S_A[3][16] = 4'hF;
    S_A[4][16] = 4'hF;
    S_A[5][16] = 4'hF;
    S_A[6][16] = 4'hF;
    S_A[7][16] = 4'hC;
    S_A[8][16] = 4'hC;
    S_A[9][16] = 4'hC;
    S_A[10][16] = 4'hC;
    S_A[11][16] = 4'hC;
    S_A[12][16] = 4'hC;
    S_A[13][16] = 4'hC;
    S_A[14][16] = 4'hC;
    S_A[15][16] = 4'hC;
    S_A[16][16] = 4'hC;
    S_A[17][16] = 4'hF;
    S_A[18][16] = 4'hF;
    S_A[19][16] = 4'hF;
    S_A[20][16] = 4'hF;
    S_A[21][16] = 4'hF;
    S_A[22][16] = 4'hF;
    S_A[23][16] = 4'hF;
    S_A[24][16] = 4'hF;
    S_A[25][16] = 4'hF;
    S_A[26][16] = 4'hF;
    S_A[27][16] = 4'hC;
    S_A[28][16] = 4'hC;
    S_A[29][16] = 4'hC;
    S_A[30][16] = 4'hC;
    S_A[31][16] = 4'hC;
    S_A[32][16] = 4'hF;
    S_A[33][16] = 4'hF;
    S_A[34][16] = 4'hF;
    S_A[35][16] = 4'hF;
    S_A[36][16] = 4'hF;
    S_A[37][16] = 4'hF;
    S_A[38][16] = 4'hF;
    S_A[39][16] = 4'hF;
    S_A[40][16] = 4'hF;
    S_A[41][16] = 4'hF;
    S_A[42][16] = 4'hF;
    S_A[43][16] = 4'hF;
    S_A[44][16] = 4'hF;
    S_A[45][16] = 4'hF;
    S_A[46][16] = 4'hF;
    S_A[47][16] = 4'hC;
    S_A[48][16] = 4'hC;
    S_A[49][16] = 4'hC;
    S_A[50][16] = 4'hC;
    S_A[51][16] = 4'hC;
    S_A[52][16] = 4'hF;
    S_A[53][16] = 4'hF;
    S_A[54][16] = 4'hF;
    S_A[55][16] = 4'hF;
    S_A[56][16] = 4'hF;
    S_A[57][16] = 4'hF;
    S_A[58][16] = 4'hF;
    S_A[59][16] = 4'hF;
    S_A[60][16] = 4'hF;
    S_A[61][16] = 4'hF;
    S_A[62][16] = 4'hC;
    S_A[63][16] = 4'hC;
    S_A[64][16] = 4'hC;
    S_A[65][16] = 4'hC;
    S_A[66][16] = 4'hC;
    S_A[67][16] = 4'hF;
    S_A[68][16] = 4'hF;
    S_A[69][16] = 4'hF;
    S_A[70][16] = 4'hF;
    S_A[71][16] = 4'hF;
    S_A[72][16] = 4'hC;
    S_A[73][16] = 4'hC;
    S_A[74][16] = 4'hC;
    S_A[75][16] = 4'hC;
    S_A[76][16] = 4'hC;
    S_A[77][16] = 4'hC;
    S_A[78][16] = 4'hC;
    S_A[79][16] = 4'hC;
    S_A[80][16] = 4'hC;
    S_A[81][16] = 4'hC;
    S_A[82][16] = 4'hF;
    S_A[83][16] = 4'hF;
    S_A[84][16] = 4'hF;
    S_A[85][16] = 4'hF;
    S_A[86][16] = 4'hF;
    S_A[87][16] = 4'hF;
    S_A[88][16] = 4'hF;
    S_A[89][16] = 4'hF;
    S_A[90][16] = 4'hF;
    S_A[91][16] = 4'hF;
    S_A[92][16] = 4'hC;
    S_A[93][16] = 4'hC;
    S_A[94][16] = 4'hC;
    S_A[95][16] = 4'hC;
    S_A[96][16] = 4'hC;
    S_A[97][16] = 4'hF;
    S_A[98][16] = 4'hF;
    S_A[99][16] = 4'hF;
    S_A[100][16] = 4'hF;
    S_A[101][16] = 4'hF;
    S_A[102][16] = 4'hC;
    S_A[103][16] = 4'hC;
    S_A[104][16] = 4'hC;
    S_A[105][16] = 4'hC;
    S_A[106][16] = 4'hC;
    S_A[107][16] = 4'hC;
    S_A[108][16] = 4'hC;
    S_A[109][16] = 4'hC;
    S_A[110][16] = 4'hC;
    S_A[111][16] = 4'hC;
    S_A[112][16] = 4'hF;
    S_A[113][16] = 4'hF;
    S_A[114][16] = 4'hF;
    S_A[0][17] = 4'hF;
    S_A[1][17] = 4'hF;
    S_A[2][17] = 4'hF;
    S_A[3][17] = 4'hF;
    S_A[4][17] = 4'hF;
    S_A[5][17] = 4'hF;
    S_A[6][17] = 4'hF;
    S_A[7][17] = 4'hF;
    S_A[8][17] = 4'hF;
    S_A[9][17] = 4'hF;
    S_A[10][17] = 4'hF;
    S_A[11][17] = 4'hF;
    S_A[12][17] = 4'hF;
    S_A[13][17] = 4'hF;
    S_A[14][17] = 4'hF;
    S_A[15][17] = 4'hF;
    S_A[16][17] = 4'hF;
    S_A[17][17] = 4'hC;
    S_A[18][17] = 4'hC;
    S_A[19][17] = 4'hC;
    S_A[20][17] = 4'hC;
    S_A[21][17] = 4'hC;
    S_A[22][17] = 4'hF;
    S_A[23][17] = 4'hF;
    S_A[24][17] = 4'hF;
    S_A[25][17] = 4'hF;
    S_A[26][17] = 4'hF;
    S_A[27][17] = 4'hC;
    S_A[28][17] = 4'hC;
    S_A[29][17] = 4'hC;
    S_A[30][17] = 4'hC;
    S_A[31][17] = 4'hC;
    S_A[32][17] = 4'hF;
    S_A[33][17] = 4'hF;
    S_A[34][17] = 4'hF;
    S_A[35][17] = 4'hF;
    S_A[36][17] = 4'hF;
    S_A[37][17] = 4'hF;
    S_A[38][17] = 4'hF;
    S_A[39][17] = 4'hF;
    S_A[40][17] = 4'hF;
    S_A[41][17] = 4'hF;
    S_A[42][17] = 4'hF;
    S_A[43][17] = 4'hF;
    S_A[44][17] = 4'hF;
    S_A[45][17] = 4'hF;
    S_A[46][17] = 4'hF;
    S_A[47][17] = 4'hC;
    S_A[48][17] = 4'hC;
    S_A[49][17] = 4'hC;
    S_A[50][17] = 4'hC;
    S_A[51][17] = 4'hC;
    S_A[52][17] = 4'hF;
    S_A[53][17] = 4'hF;
    S_A[54][17] = 4'hF;
    S_A[55][17] = 4'hF;
    S_A[56][17] = 4'hF;
    S_A[57][17] = 4'hF;
    S_A[58][17] = 4'hF;
    S_A[59][17] = 4'hF;
    S_A[60][17] = 4'hF;
    S_A[61][17] = 4'hF;
    S_A[62][17] = 4'hC;
    S_A[63][17] = 4'hC;
    S_A[64][17] = 4'hC;
    S_A[65][17] = 4'hC;
    S_A[66][17] = 4'hC;
    S_A[67][17] = 4'hF;
    S_A[68][17] = 4'hF;
    S_A[69][17] = 4'hF;
    S_A[70][17] = 4'hF;
    S_A[71][17] = 4'hF;
    S_A[72][17] = 4'hC;
    S_A[73][17] = 4'hC;
    S_A[74][17] = 4'hC;
    S_A[75][17] = 4'hC;
    S_A[76][17] = 4'hC;
    S_A[77][17] = 4'hF;
    S_A[78][17] = 4'hF;
    S_A[79][17] = 4'hF;
    S_A[80][17] = 4'hF;
    S_A[81][17] = 4'hF;
    S_A[82][17] = 4'hF;
    S_A[83][17] = 4'hF;
    S_A[84][17] = 4'hF;
    S_A[85][17] = 4'hF;
    S_A[86][17] = 4'hF;
    S_A[87][17] = 4'hF;
    S_A[88][17] = 4'hF;
    S_A[89][17] = 4'hF;
    S_A[90][17] = 4'hF;
    S_A[91][17] = 4'hF;
    S_A[92][17] = 4'hC;
    S_A[93][17] = 4'hC;
    S_A[94][17] = 4'hC;
    S_A[95][17] = 4'hC;
    S_A[96][17] = 4'hC;
    S_A[97][17] = 4'hC;
    S_A[98][17] = 4'hC;
    S_A[99][17] = 4'hC;
    S_A[100][17] = 4'hC;
    S_A[101][17] = 4'hC;
    S_A[102][17] = 4'hF;
    S_A[103][17] = 4'hF;
    S_A[104][17] = 4'hF;
    S_A[105][17] = 4'hF;
    S_A[106][17] = 4'hF;
    S_A[107][17] = 4'hF;
    S_A[108][17] = 4'hF;
    S_A[109][17] = 4'hF;
    S_A[110][17] = 4'hF;
    S_A[111][17] = 4'hF;
    S_A[112][17] = 4'hF;
    S_A[113][17] = 4'hF;
    S_A[114][17] = 4'hF;
    S_A[0][18] = 4'hF;
    S_A[1][18] = 4'hF;
    S_A[2][18] = 4'hF;
    S_A[3][18] = 4'hF;
    S_A[4][18] = 4'hF;
    S_A[5][18] = 4'hF;
    S_A[6][18] = 4'hF;
    S_A[7][18] = 4'hF;
    S_A[8][18] = 4'hF;
    S_A[9][18] = 4'hF;
    S_A[10][18] = 4'hF;
    S_A[11][18] = 4'hF;
    S_A[12][18] = 4'hF;
    S_A[13][18] = 4'hF;
    S_A[14][18] = 4'hF;
    S_A[15][18] = 4'hF;
    S_A[16][18] = 4'hF;
    S_A[17][18] = 4'hC;
    S_A[18][18] = 4'hC;
    S_A[19][18] = 4'hC;
    S_A[20][18] = 4'hC;
    S_A[21][18] = 4'hC;
    S_A[22][18] = 4'hF;
    S_A[23][18] = 4'hF;
    S_A[24][18] = 4'hF;
    S_A[25][18] = 4'hF;
    S_A[26][18] = 4'hF;
    S_A[27][18] = 4'hC;
    S_A[28][18] = 4'hC;
    S_A[29][18] = 4'hC;
    S_A[30][18] = 4'hC;
    S_A[31][18] = 4'hC;
    S_A[32][18] = 4'hF;
    S_A[33][18] = 4'hF;
    S_A[34][18] = 4'hF;
    S_A[35][18] = 4'hF;
    S_A[36][18] = 4'hF;
    S_A[37][18] = 4'hF;
    S_A[38][18] = 4'hF;
    S_A[39][18] = 4'hF;
    S_A[40][18] = 4'hF;
    S_A[41][18] = 4'hF;
    S_A[42][18] = 4'hF;
    S_A[43][18] = 4'hF;
    S_A[44][18] = 4'hF;
    S_A[45][18] = 4'hF;
    S_A[46][18] = 4'hF;
    S_A[47][18] = 4'hC;
    S_A[48][18] = 4'hC;
    S_A[49][18] = 4'hC;
    S_A[50][18] = 4'hC;
    S_A[51][18] = 4'hC;
    S_A[52][18] = 4'hF;
    S_A[53][18] = 4'hF;
    S_A[54][18] = 4'hF;
    S_A[55][18] = 4'hF;
    S_A[56][18] = 4'hF;
    S_A[57][18] = 4'hF;
    S_A[58][18] = 4'hF;
    S_A[59][18] = 4'hF;
    S_A[60][18] = 4'hF;
    S_A[61][18] = 4'hF;
    S_A[62][18] = 4'hC;
    S_A[63][18] = 4'hC;
    S_A[64][18] = 4'hC;
    S_A[65][18] = 4'hC;
    S_A[66][18] = 4'hC;
    S_A[67][18] = 4'hF;
    S_A[68][18] = 4'hF;
    S_A[69][18] = 4'hF;
    S_A[70][18] = 4'hF;
    S_A[71][18] = 4'hF;
    S_A[72][18] = 4'hC;
    S_A[73][18] = 4'hC;
    S_A[74][18] = 4'hC;
    S_A[75][18] = 4'hC;
    S_A[76][18] = 4'hC;
    S_A[77][18] = 4'hF;
    S_A[78][18] = 4'hF;
    S_A[79][18] = 4'hF;
    S_A[80][18] = 4'hF;
    S_A[81][18] = 4'hF;
    S_A[82][18] = 4'hF;
    S_A[83][18] = 4'hF;
    S_A[84][18] = 4'hF;
    S_A[85][18] = 4'hF;
    S_A[86][18] = 4'hF;
    S_A[87][18] = 4'hF;
    S_A[88][18] = 4'hF;
    S_A[89][18] = 4'hF;
    S_A[90][18] = 4'hF;
    S_A[91][18] = 4'hF;
    S_A[92][18] = 4'hC;
    S_A[93][18] = 4'hC;
    S_A[94][18] = 4'hC;
    S_A[95][18] = 4'hC;
    S_A[96][18] = 4'hC;
    S_A[97][18] = 4'hC;
    S_A[98][18] = 4'hC;
    S_A[99][18] = 4'hC;
    S_A[100][18] = 4'hC;
    S_A[101][18] = 4'hC;
    S_A[102][18] = 4'hF;
    S_A[103][18] = 4'hF;
    S_A[104][18] = 4'hF;
    S_A[105][18] = 4'hF;
    S_A[106][18] = 4'hF;
    S_A[107][18] = 4'hF;
    S_A[108][18] = 4'hF;
    S_A[109][18] = 4'hF;
    S_A[110][18] = 4'hF;
    S_A[111][18] = 4'hF;
    S_A[112][18] = 4'hF;
    S_A[113][18] = 4'hF;
    S_A[114][18] = 4'hF;
    S_A[0][19] = 4'hF;
    S_A[1][19] = 4'hF;
    S_A[2][19] = 4'hF;
    S_A[3][19] = 4'hF;
    S_A[4][19] = 4'hF;
    S_A[5][19] = 4'hF;
    S_A[6][19] = 4'hF;
    S_A[7][19] = 4'hF;
    S_A[8][19] = 4'hF;
    S_A[9][19] = 4'hF;
    S_A[10][19] = 4'hF;
    S_A[11][19] = 4'hF;
    S_A[12][19] = 4'hF;
    S_A[13][19] = 4'hF;
    S_A[14][19] = 4'hF;
    S_A[15][19] = 4'hF;
    S_A[16][19] = 4'hF;
    S_A[17][19] = 4'hC;
    S_A[18][19] = 4'hC;
    S_A[19][19] = 4'hC;
    S_A[20][19] = 4'hC;
    S_A[21][19] = 4'hC;
    S_A[22][19] = 4'hF;
    S_A[23][19] = 4'hF;
    S_A[24][19] = 4'hF;
    S_A[25][19] = 4'hF;
    S_A[26][19] = 4'hF;
    S_A[27][19] = 4'hC;
    S_A[28][19] = 4'hC;
    S_A[29][19] = 4'hC;
    S_A[30][19] = 4'hC;
    S_A[31][19] = 4'hC;
    S_A[32][19] = 4'hF;
    S_A[33][19] = 4'hF;
    S_A[34][19] = 4'hF;
    S_A[35][19] = 4'hF;
    S_A[36][19] = 4'hF;
    S_A[37][19] = 4'hF;
    S_A[38][19] = 4'hF;
    S_A[39][19] = 4'hF;
    S_A[40][19] = 4'hF;
    S_A[41][19] = 4'hF;
    S_A[42][19] = 4'hF;
    S_A[43][19] = 4'hF;
    S_A[44][19] = 4'hF;
    S_A[45][19] = 4'hF;
    S_A[46][19] = 4'hF;
    S_A[47][19] = 4'hC;
    S_A[48][19] = 4'hC;
    S_A[49][19] = 4'hC;
    S_A[50][19] = 4'hC;
    S_A[51][19] = 4'hC;
    S_A[52][19] = 4'hF;
    S_A[53][19] = 4'hF;
    S_A[54][19] = 4'hF;
    S_A[55][19] = 4'hF;
    S_A[56][19] = 4'hF;
    S_A[57][19] = 4'hF;
    S_A[58][19] = 4'hF;
    S_A[59][19] = 4'hF;
    S_A[60][19] = 4'hF;
    S_A[61][19] = 4'hF;
    S_A[62][19] = 4'hC;
    S_A[63][19] = 4'hC;
    S_A[64][19] = 4'hC;
    S_A[65][19] = 4'hC;
    S_A[66][19] = 4'hC;
    S_A[67][19] = 4'hF;
    S_A[68][19] = 4'hF;
    S_A[69][19] = 4'hF;
    S_A[70][19] = 4'hF;
    S_A[71][19] = 4'hF;
    S_A[72][19] = 4'hC;
    S_A[73][19] = 4'hC;
    S_A[74][19] = 4'hC;
    S_A[75][19] = 4'hC;
    S_A[76][19] = 4'hC;
    S_A[77][19] = 4'hF;
    S_A[78][19] = 4'hF;
    S_A[79][19] = 4'hF;
    S_A[80][19] = 4'hF;
    S_A[81][19] = 4'hF;
    S_A[82][19] = 4'hF;
    S_A[83][19] = 4'hF;
    S_A[84][19] = 4'hF;
    S_A[85][19] = 4'hF;
    S_A[86][19] = 4'hF;
    S_A[87][19] = 4'hF;
    S_A[88][19] = 4'hF;
    S_A[89][19] = 4'hF;
    S_A[90][19] = 4'hF;
    S_A[91][19] = 4'hF;
    S_A[92][19] = 4'hC;
    S_A[93][19] = 4'hC;
    S_A[94][19] = 4'hC;
    S_A[95][19] = 4'hC;
    S_A[96][19] = 4'hC;
    S_A[97][19] = 4'hC;
    S_A[98][19] = 4'hC;
    S_A[99][19] = 4'hC;
    S_A[100][19] = 4'hC;
    S_A[101][19] = 4'hC;
    S_A[102][19] = 4'hF;
    S_A[103][19] = 4'hF;
    S_A[104][19] = 4'hF;
    S_A[105][19] = 4'hF;
    S_A[106][19] = 4'hF;
    S_A[107][19] = 4'hF;
    S_A[108][19] = 4'hF;
    S_A[109][19] = 4'hF;
    S_A[110][19] = 4'hF;
    S_A[111][19] = 4'hF;
    S_A[112][19] = 4'hF;
    S_A[113][19] = 4'hF;
    S_A[114][19] = 4'hF;
    S_A[0][20] = 4'hF;
    S_A[1][20] = 4'hF;
    S_A[2][20] = 4'hF;
    S_A[3][20] = 4'hF;
    S_A[4][20] = 4'hF;
    S_A[5][20] = 4'hF;
    S_A[6][20] = 4'hF;
    S_A[7][20] = 4'hF;
    S_A[8][20] = 4'hF;
    S_A[9][20] = 4'hF;
    S_A[10][20] = 4'hF;
    S_A[11][20] = 4'hF;
    S_A[12][20] = 4'hF;
    S_A[13][20] = 4'hF;
    S_A[14][20] = 4'hF;
    S_A[15][20] = 4'hF;
    S_A[16][20] = 4'hF;
    S_A[17][20] = 4'hC;
    S_A[18][20] = 4'hC;
    S_A[19][20] = 4'hC;
    S_A[20][20] = 4'hC;
    S_A[21][20] = 4'hC;
    S_A[22][20] = 4'hF;
    S_A[23][20] = 4'hF;
    S_A[24][20] = 4'hF;
    S_A[25][20] = 4'hF;
    S_A[26][20] = 4'hF;
    S_A[27][20] = 4'hC;
    S_A[28][20] = 4'hC;
    S_A[29][20] = 4'hC;
    S_A[30][20] = 4'hC;
    S_A[31][20] = 4'hC;
    S_A[32][20] = 4'hF;
    S_A[33][20] = 4'hF;
    S_A[34][20] = 4'hF;
    S_A[35][20] = 4'hF;
    S_A[36][20] = 4'hF;
    S_A[37][20] = 4'hF;
    S_A[38][20] = 4'hF;
    S_A[39][20] = 4'hF;
    S_A[40][20] = 4'hF;
    S_A[41][20] = 4'hF;
    S_A[42][20] = 4'hF;
    S_A[43][20] = 4'hF;
    S_A[44][20] = 4'hF;
    S_A[45][20] = 4'hF;
    S_A[46][20] = 4'hF;
    S_A[47][20] = 4'hC;
    S_A[48][20] = 4'hC;
    S_A[49][20] = 4'hC;
    S_A[50][20] = 4'hC;
    S_A[51][20] = 4'hC;
    S_A[52][20] = 4'hF;
    S_A[53][20] = 4'hF;
    S_A[54][20] = 4'hF;
    S_A[55][20] = 4'hF;
    S_A[56][20] = 4'hF;
    S_A[57][20] = 4'hF;
    S_A[58][20] = 4'hF;
    S_A[59][20] = 4'hF;
    S_A[60][20] = 4'hF;
    S_A[61][20] = 4'hF;
    S_A[62][20] = 4'hC;
    S_A[63][20] = 4'hC;
    S_A[64][20] = 4'hC;
    S_A[65][20] = 4'hC;
    S_A[66][20] = 4'hC;
    S_A[67][20] = 4'hF;
    S_A[68][20] = 4'hF;
    S_A[69][20] = 4'hF;
    S_A[70][20] = 4'hF;
    S_A[71][20] = 4'hF;
    S_A[72][20] = 4'hC;
    S_A[73][20] = 4'hC;
    S_A[74][20] = 4'hC;
    S_A[75][20] = 4'hC;
    S_A[76][20] = 4'hC;
    S_A[77][20] = 4'hF;
    S_A[78][20] = 4'hF;
    S_A[79][20] = 4'hF;
    S_A[80][20] = 4'hF;
    S_A[81][20] = 4'hF;
    S_A[82][20] = 4'hF;
    S_A[83][20] = 4'hF;
    S_A[84][20] = 4'hF;
    S_A[85][20] = 4'hF;
    S_A[86][20] = 4'hF;
    S_A[87][20] = 4'hF;
    S_A[88][20] = 4'hF;
    S_A[89][20] = 4'hF;
    S_A[90][20] = 4'hF;
    S_A[91][20] = 4'hF;
    S_A[92][20] = 4'hC;
    S_A[93][20] = 4'hC;
    S_A[94][20] = 4'hC;
    S_A[95][20] = 4'hC;
    S_A[96][20] = 4'hC;
    S_A[97][20] = 4'hC;
    S_A[98][20] = 4'hC;
    S_A[99][20] = 4'hC;
    S_A[100][20] = 4'hC;
    S_A[101][20] = 4'hC;
    S_A[102][20] = 4'hF;
    S_A[103][20] = 4'hF;
    S_A[104][20] = 4'hF;
    S_A[105][20] = 4'hF;
    S_A[106][20] = 4'hF;
    S_A[107][20] = 4'hF;
    S_A[108][20] = 4'hF;
    S_A[109][20] = 4'hF;
    S_A[110][20] = 4'hF;
    S_A[111][20] = 4'hF;
    S_A[112][20] = 4'hF;
    S_A[113][20] = 4'hF;
    S_A[114][20] = 4'hF;
    S_A[0][21] = 4'hF;
    S_A[1][21] = 4'hF;
    S_A[2][21] = 4'hF;
    S_A[3][21] = 4'hF;
    S_A[4][21] = 4'hF;
    S_A[5][21] = 4'hF;
    S_A[6][21] = 4'hF;
    S_A[7][21] = 4'hF;
    S_A[8][21] = 4'hF;
    S_A[9][21] = 4'hF;
    S_A[10][21] = 4'hF;
    S_A[11][21] = 4'hF;
    S_A[12][21] = 4'hF;
    S_A[13][21] = 4'hF;
    S_A[14][21] = 4'hF;
    S_A[15][21] = 4'hF;
    S_A[16][21] = 4'hF;
    S_A[17][21] = 4'hC;
    S_A[18][21] = 4'hC;
    S_A[19][21] = 4'hC;
    S_A[20][21] = 4'hC;
    S_A[21][21] = 4'hC;
    S_A[22][21] = 4'hF;
    S_A[23][21] = 4'hF;
    S_A[24][21] = 4'hF;
    S_A[25][21] = 4'hF;
    S_A[26][21] = 4'hF;
    S_A[27][21] = 4'hC;
    S_A[28][21] = 4'hC;
    S_A[29][21] = 4'hC;
    S_A[30][21] = 4'hC;
    S_A[31][21] = 4'hC;
    S_A[32][21] = 4'hF;
    S_A[33][21] = 4'hF;
    S_A[34][21] = 4'hF;
    S_A[35][21] = 4'hF;
    S_A[36][21] = 4'hF;
    S_A[37][21] = 4'hF;
    S_A[38][21] = 4'hF;
    S_A[39][21] = 4'hF;
    S_A[40][21] = 4'hF;
    S_A[41][21] = 4'hF;
    S_A[42][21] = 4'hF;
    S_A[43][21] = 4'hF;
    S_A[44][21] = 4'hF;
    S_A[45][21] = 4'hF;
    S_A[46][21] = 4'hF;
    S_A[47][21] = 4'hC;
    S_A[48][21] = 4'hC;
    S_A[49][21] = 4'hC;
    S_A[50][21] = 4'hC;
    S_A[51][21] = 4'hC;
    S_A[52][21] = 4'hF;
    S_A[53][21] = 4'hF;
    S_A[54][21] = 4'hF;
    S_A[55][21] = 4'hF;
    S_A[56][21] = 4'hF;
    S_A[57][21] = 4'hF;
    S_A[58][21] = 4'hF;
    S_A[59][21] = 4'hF;
    S_A[60][21] = 4'hF;
    S_A[61][21] = 4'hF;
    S_A[62][21] = 4'hC;
    S_A[63][21] = 4'hC;
    S_A[64][21] = 4'hC;
    S_A[65][21] = 4'hC;
    S_A[66][21] = 4'hC;
    S_A[67][21] = 4'hF;
    S_A[68][21] = 4'hF;
    S_A[69][21] = 4'hF;
    S_A[70][21] = 4'hF;
    S_A[71][21] = 4'hF;
    S_A[72][21] = 4'hC;
    S_A[73][21] = 4'hC;
    S_A[74][21] = 4'hC;
    S_A[75][21] = 4'hC;
    S_A[76][21] = 4'hC;
    S_A[77][21] = 4'hF;
    S_A[78][21] = 4'hF;
    S_A[79][21] = 4'hF;
    S_A[80][21] = 4'hF;
    S_A[81][21] = 4'hF;
    S_A[82][21] = 4'hF;
    S_A[83][21] = 4'hF;
    S_A[84][21] = 4'hF;
    S_A[85][21] = 4'hF;
    S_A[86][21] = 4'hF;
    S_A[87][21] = 4'hF;
    S_A[88][21] = 4'hF;
    S_A[89][21] = 4'hF;
    S_A[90][21] = 4'hF;
    S_A[91][21] = 4'hF;
    S_A[92][21] = 4'hC;
    S_A[93][21] = 4'hC;
    S_A[94][21] = 4'hC;
    S_A[95][21] = 4'hC;
    S_A[96][21] = 4'hC;
    S_A[97][21] = 4'hC;
    S_A[98][21] = 4'hC;
    S_A[99][21] = 4'hC;
    S_A[100][21] = 4'hC;
    S_A[101][21] = 4'hC;
    S_A[102][21] = 4'hF;
    S_A[103][21] = 4'hF;
    S_A[104][21] = 4'hF;
    S_A[105][21] = 4'hF;
    S_A[106][21] = 4'hF;
    S_A[107][21] = 4'hF;
    S_A[108][21] = 4'hF;
    S_A[109][21] = 4'hF;
    S_A[110][21] = 4'hF;
    S_A[111][21] = 4'hF;
    S_A[112][21] = 4'hF;
    S_A[113][21] = 4'hF;
    S_A[114][21] = 4'hF;
    S_A[0][22] = 4'hF;
    S_A[1][22] = 4'hF;
    S_A[2][22] = 4'hC;
    S_A[3][22] = 4'hC;
    S_A[4][22] = 4'hC;
    S_A[5][22] = 4'hC;
    S_A[6][22] = 4'hC;
    S_A[7][22] = 4'hC;
    S_A[8][22] = 4'hC;
    S_A[9][22] = 4'hC;
    S_A[10][22] = 4'hC;
    S_A[11][22] = 4'hC;
    S_A[12][22] = 4'hC;
    S_A[13][22] = 4'hC;
    S_A[14][22] = 4'hC;
    S_A[15][22] = 4'hC;
    S_A[16][22] = 4'hC;
    S_A[17][22] = 4'hF;
    S_A[18][22] = 4'hF;
    S_A[19][22] = 4'hF;
    S_A[20][22] = 4'hF;
    S_A[21][22] = 4'hF;
    S_A[22][22] = 4'hF;
    S_A[23][22] = 4'hF;
    S_A[24][22] = 4'hF;
    S_A[25][22] = 4'hF;
    S_A[26][22] = 4'hF;
    S_A[27][22] = 4'hF;
    S_A[28][22] = 4'hF;
    S_A[29][22] = 4'hF;
    S_A[30][22] = 4'hF;
    S_A[31][22] = 4'hF;
    S_A[32][22] = 4'hC;
    S_A[33][22] = 4'hC;
    S_A[34][22] = 4'hC;
    S_A[35][22] = 4'hC;
    S_A[36][22] = 4'hC;
    S_A[37][22] = 4'hC;
    S_A[38][22] = 4'hC;
    S_A[39][22] = 4'hC;
    S_A[40][22] = 4'hC;
    S_A[41][22] = 4'hC;
    S_A[42][22] = 4'hF;
    S_A[43][22] = 4'hF;
    S_A[44][22] = 4'hF;
    S_A[45][22] = 4'hF;
    S_A[46][22] = 4'hF;
    S_A[47][22] = 4'hF;
    S_A[48][22] = 4'hF;
    S_A[49][22] = 4'hF;
    S_A[50][22] = 4'hF;
    S_A[51][22] = 4'hF;
    S_A[52][22] = 4'hC;
    S_A[53][22] = 4'hC;
    S_A[54][22] = 4'hC;
    S_A[55][22] = 4'hC;
    S_A[56][22] = 4'hC;
    S_A[57][22] = 4'hC;
    S_A[58][22] = 4'hC;
    S_A[59][22] = 4'hC;
    S_A[60][22] = 4'hC;
    S_A[61][22] = 4'hC;
    S_A[62][22] = 4'hF;
    S_A[63][22] = 4'hF;
    S_A[64][22] = 4'hF;
    S_A[65][22] = 4'hF;
    S_A[66][22] = 4'hF;
    S_A[67][22] = 4'hF;
    S_A[68][22] = 4'hF;
    S_A[69][22] = 4'hF;
    S_A[70][22] = 4'hF;
    S_A[71][22] = 4'hF;
    S_A[72][22] = 4'hC;
    S_A[73][22] = 4'hC;
    S_A[74][22] = 4'hC;
    S_A[75][22] = 4'hC;
    S_A[76][22] = 4'hC;
    S_A[77][22] = 4'hF;
    S_A[78][22] = 4'hF;
    S_A[79][22] = 4'hF;
    S_A[80][22] = 4'hF;
    S_A[81][22] = 4'hF;
    S_A[82][22] = 4'hF;
    S_A[83][22] = 4'hF;
    S_A[84][22] = 4'hF;
    S_A[85][22] = 4'hF;
    S_A[86][22] = 4'hF;
    S_A[87][22] = 4'hF;
    S_A[88][22] = 4'hF;
    S_A[89][22] = 4'hF;
    S_A[90][22] = 4'hF;
    S_A[91][22] = 4'hF;
    S_A[92][22] = 4'hF;
    S_A[93][22] = 4'hF;
    S_A[94][22] = 4'hF;
    S_A[95][22] = 4'hF;
    S_A[96][22] = 4'hF;
    S_A[97][22] = 4'hC;
    S_A[98][22] = 4'hC;
    S_A[99][22] = 4'hC;
    S_A[100][22] = 4'hC;
    S_A[101][22] = 4'hC;
    S_A[102][22] = 4'hC;
    S_A[103][22] = 4'hC;
    S_A[104][22] = 4'hC;
    S_A[105][22] = 4'hC;
    S_A[106][22] = 4'hC;
    S_A[107][22] = 4'hF;
    S_A[108][22] = 4'hF;
    S_A[109][22] = 4'hF;
    S_A[110][22] = 4'hF;
    S_A[111][22] = 4'hF;
    S_A[112][22] = 4'hF;
    S_A[113][22] = 4'hF;
    S_A[114][22] = 4'hF;
    S_A[0][23] = 4'hF;
    S_A[1][23] = 4'hF;
    S_A[2][23] = 4'hC;
    S_A[3][23] = 4'hC;
    S_A[4][23] = 4'hC;
    S_A[5][23] = 4'hC;
    S_A[6][23] = 4'hC;
    S_A[7][23] = 4'hC;
    S_A[8][23] = 4'hC;
    S_A[9][23] = 4'hC;
    S_A[10][23] = 4'hC;
    S_A[11][23] = 4'hC;
    S_A[12][23] = 4'hC;
    S_A[13][23] = 4'hC;
    S_A[14][23] = 4'hC;
    S_A[15][23] = 4'hC;
    S_A[16][23] = 4'hC;
    S_A[17][23] = 4'hF;
    S_A[18][23] = 4'hF;
    S_A[19][23] = 4'hF;
    S_A[20][23] = 4'hF;
    S_A[21][23] = 4'hF;
    S_A[22][23] = 4'hF;
    S_A[23][23] = 4'hF;
    S_A[24][23] = 4'hF;
    S_A[25][23] = 4'hF;
    S_A[26][23] = 4'hF;
    S_A[27][23] = 4'hF;
    S_A[28][23] = 4'hF;
    S_A[29][23] = 4'hF;
    S_A[30][23] = 4'hF;
    S_A[31][23] = 4'hF;
    S_A[32][23] = 4'hC;
    S_A[33][23] = 4'hC;
    S_A[34][23] = 4'hC;
    S_A[35][23] = 4'hC;
    S_A[36][23] = 4'hC;
    S_A[37][23] = 4'hC;
    S_A[38][23] = 4'hC;
    S_A[39][23] = 4'hC;
    S_A[40][23] = 4'hC;
    S_A[41][23] = 4'hC;
    S_A[42][23] = 4'hF;
    S_A[43][23] = 4'hF;
    S_A[44][23] = 4'hF;
    S_A[45][23] = 4'hF;
    S_A[46][23] = 4'hF;
    S_A[47][23] = 4'hF;
    S_A[48][23] = 4'hF;
    S_A[49][23] = 4'hF;
    S_A[50][23] = 4'hF;
    S_A[51][23] = 4'hF;
    S_A[52][23] = 4'hC;
    S_A[53][23] = 4'hC;
    S_A[54][23] = 4'hC;
    S_A[55][23] = 4'hC;
    S_A[56][23] = 4'hC;
    S_A[57][23] = 4'hC;
    S_A[58][23] = 4'hC;
    S_A[59][23] = 4'hC;
    S_A[60][23] = 4'hC;
    S_A[61][23] = 4'hC;
    S_A[62][23] = 4'hF;
    S_A[63][23] = 4'hF;
    S_A[64][23] = 4'hF;
    S_A[65][23] = 4'hF;
    S_A[66][23] = 4'hF;
    S_A[67][23] = 4'hF;
    S_A[68][23] = 4'hF;
    S_A[69][23] = 4'hF;
    S_A[70][23] = 4'hF;
    S_A[71][23] = 4'hF;
    S_A[72][23] = 4'hC;
    S_A[73][23] = 4'hC;
    S_A[74][23] = 4'hC;
    S_A[75][23] = 4'hC;
    S_A[76][23] = 4'hC;
    S_A[77][23] = 4'hF;
    S_A[78][23] = 4'hF;
    S_A[79][23] = 4'hF;
    S_A[80][23] = 4'hF;
    S_A[81][23] = 4'hF;
    S_A[82][23] = 4'hF;
    S_A[83][23] = 4'hF;
    S_A[84][23] = 4'hF;
    S_A[85][23] = 4'hF;
    S_A[86][23] = 4'hF;
    S_A[87][23] = 4'hF;
    S_A[88][23] = 4'hF;
    S_A[89][23] = 4'hF;
    S_A[90][23] = 4'hF;
    S_A[91][23] = 4'hF;
    S_A[92][23] = 4'hF;
    S_A[93][23] = 4'hF;
    S_A[94][23] = 4'hF;
    S_A[95][23] = 4'hF;
    S_A[96][23] = 4'hF;
    S_A[97][23] = 4'hC;
    S_A[98][23] = 4'hC;
    S_A[99][23] = 4'hC;
    S_A[100][23] = 4'hC;
    S_A[101][23] = 4'hC;
    S_A[102][23] = 4'hC;
    S_A[103][23] = 4'hC;
    S_A[104][23] = 4'hC;
    S_A[105][23] = 4'hC;
    S_A[106][23] = 4'hC;
    S_A[107][23] = 4'hF;
    S_A[108][23] = 4'hF;
    S_A[109][23] = 4'hF;
    S_A[110][23] = 4'hF;
    S_A[111][23] = 4'hF;
    S_A[112][23] = 4'hF;
    S_A[113][23] = 4'hF;
    S_A[114][23] = 4'hF;
    S_A[0][24] = 4'hF;
    S_A[1][24] = 4'hF;
    S_A[2][24] = 4'hC;
    S_A[3][24] = 4'hC;
    S_A[4][24] = 4'hC;
    S_A[5][24] = 4'hC;
    S_A[6][24] = 4'hC;
    S_A[7][24] = 4'hC;
    S_A[8][24] = 4'hC;
    S_A[9][24] = 4'hC;
    S_A[10][24] = 4'hC;
    S_A[11][24] = 4'hC;
    S_A[12][24] = 4'hC;
    S_A[13][24] = 4'hC;
    S_A[14][24] = 4'hC;
    S_A[15][24] = 4'hC;
    S_A[16][24] = 4'hC;
    S_A[17][24] = 4'hF;
    S_A[18][24] = 4'hF;
    S_A[19][24] = 4'hF;
    S_A[20][24] = 4'hF;
    S_A[21][24] = 4'hF;
    S_A[22][24] = 4'hF;
    S_A[23][24] = 4'hF;
    S_A[24][24] = 4'hF;
    S_A[25][24] = 4'hF;
    S_A[26][24] = 4'hF;
    S_A[27][24] = 4'hF;
    S_A[28][24] = 4'hF;
    S_A[29][24] = 4'hF;
    S_A[30][24] = 4'hF;
    S_A[31][24] = 4'hF;
    S_A[32][24] = 4'hC;
    S_A[33][24] = 4'hC;
    S_A[34][24] = 4'hC;
    S_A[35][24] = 4'hC;
    S_A[36][24] = 4'hC;
    S_A[37][24] = 4'hC;
    S_A[38][24] = 4'hC;
    S_A[39][24] = 4'hC;
    S_A[40][24] = 4'hC;
    S_A[41][24] = 4'hC;
    S_A[42][24] = 4'hF;
    S_A[43][24] = 4'hF;
    S_A[44][24] = 4'hF;
    S_A[45][24] = 4'hF;
    S_A[46][24] = 4'hF;
    S_A[47][24] = 4'hF;
    S_A[48][24] = 4'hF;
    S_A[49][24] = 4'hF;
    S_A[50][24] = 4'hF;
    S_A[51][24] = 4'hF;
    S_A[52][24] = 4'hC;
    S_A[53][24] = 4'hC;
    S_A[54][24] = 4'hC;
    S_A[55][24] = 4'hC;
    S_A[56][24] = 4'hC;
    S_A[57][24] = 4'hC;
    S_A[58][24] = 4'hC;
    S_A[59][24] = 4'hC;
    S_A[60][24] = 4'hC;
    S_A[61][24] = 4'hC;
    S_A[62][24] = 4'hF;
    S_A[63][24] = 4'hF;
    S_A[64][24] = 4'hF;
    S_A[65][24] = 4'hF;
    S_A[66][24] = 4'hF;
    S_A[67][24] = 4'hF;
    S_A[68][24] = 4'hF;
    S_A[69][24] = 4'hF;
    S_A[70][24] = 4'hF;
    S_A[71][24] = 4'hF;
    S_A[72][24] = 4'hC;
    S_A[73][24] = 4'hC;
    S_A[74][24] = 4'hC;
    S_A[75][24] = 4'hC;
    S_A[76][24] = 4'hC;
    S_A[77][24] = 4'hF;
    S_A[78][24] = 4'hF;
    S_A[79][24] = 4'hF;
    S_A[80][24] = 4'hF;
    S_A[81][24] = 4'hF;
    S_A[82][24] = 4'hF;
    S_A[83][24] = 4'hF;
    S_A[84][24] = 4'hF;
    S_A[85][24] = 4'hF;
    S_A[86][24] = 4'hF;
    S_A[87][24] = 4'hF;
    S_A[88][24] = 4'hF;
    S_A[89][24] = 4'hF;
    S_A[90][24] = 4'hF;
    S_A[91][24] = 4'hF;
    S_A[92][24] = 4'hF;
    S_A[93][24] = 4'hF;
    S_A[94][24] = 4'hF;
    S_A[95][24] = 4'hF;
    S_A[96][24] = 4'hF;
    S_A[97][24] = 4'hC;
    S_A[98][24] = 4'hC;
    S_A[99][24] = 4'hC;
    S_A[100][24] = 4'hC;
    S_A[101][24] = 4'hC;
    S_A[102][24] = 4'hC;
    S_A[103][24] = 4'hC;
    S_A[104][24] = 4'hC;
    S_A[105][24] = 4'hC;
    S_A[106][24] = 4'hC;
    S_A[107][24] = 4'hF;
    S_A[108][24] = 4'hF;
    S_A[109][24] = 4'hF;
    S_A[110][24] = 4'hF;
    S_A[111][24] = 4'hF;
    S_A[112][24] = 4'hF;
    S_A[113][24] = 4'hF;
    S_A[114][24] = 4'hF;
    S_A[0][25] = 4'hF;
    S_A[1][25] = 4'hF;
    S_A[2][25] = 4'hC;
    S_A[3][25] = 4'hC;
    S_A[4][25] = 4'hC;
    S_A[5][25] = 4'hC;
    S_A[6][25] = 4'hC;
    S_A[7][25] = 4'hC;
    S_A[8][25] = 4'hC;
    S_A[9][25] = 4'hC;
    S_A[10][25] = 4'hC;
    S_A[11][25] = 4'hC;
    S_A[12][25] = 4'hC;
    S_A[13][25] = 4'hC;
    S_A[14][25] = 4'hC;
    S_A[15][25] = 4'hC;
    S_A[16][25] = 4'hC;
    S_A[17][25] = 4'hF;
    S_A[18][25] = 4'hF;
    S_A[19][25] = 4'hF;
    S_A[20][25] = 4'hF;
    S_A[21][25] = 4'hF;
    S_A[22][25] = 4'hF;
    S_A[23][25] = 4'hF;
    S_A[24][25] = 4'hF;
    S_A[25][25] = 4'hF;
    S_A[26][25] = 4'hF;
    S_A[27][25] = 4'hF;
    S_A[28][25] = 4'hF;
    S_A[29][25] = 4'hF;
    S_A[30][25] = 4'hF;
    S_A[31][25] = 4'hF;
    S_A[32][25] = 4'hC;
    S_A[33][25] = 4'hC;
    S_A[34][25] = 4'hC;
    S_A[35][25] = 4'hC;
    S_A[36][25] = 4'hC;
    S_A[37][25] = 4'hC;
    S_A[38][25] = 4'hC;
    S_A[39][25] = 4'hC;
    S_A[40][25] = 4'hC;
    S_A[41][25] = 4'hC;
    S_A[42][25] = 4'hF;
    S_A[43][25] = 4'hF;
    S_A[44][25] = 4'hF;
    S_A[45][25] = 4'hF;
    S_A[46][25] = 4'hF;
    S_A[47][25] = 4'hF;
    S_A[48][25] = 4'hF;
    S_A[49][25] = 4'hF;
    S_A[50][25] = 4'hF;
    S_A[51][25] = 4'hF;
    S_A[52][25] = 4'hC;
    S_A[53][25] = 4'hC;
    S_A[54][25] = 4'hC;
    S_A[55][25] = 4'hC;
    S_A[56][25] = 4'hC;
    S_A[57][25] = 4'hC;
    S_A[58][25] = 4'hC;
    S_A[59][25] = 4'hC;
    S_A[60][25] = 4'hC;
    S_A[61][25] = 4'hC;
    S_A[62][25] = 4'hF;
    S_A[63][25] = 4'hF;
    S_A[64][25] = 4'hF;
    S_A[65][25] = 4'hF;
    S_A[66][25] = 4'hF;
    S_A[67][25] = 4'hF;
    S_A[68][25] = 4'hF;
    S_A[69][25] = 4'hF;
    S_A[70][25] = 4'hF;
    S_A[71][25] = 4'hF;
    S_A[72][25] = 4'hC;
    S_A[73][25] = 4'hC;
    S_A[74][25] = 4'hC;
    S_A[75][25] = 4'hC;
    S_A[76][25] = 4'hC;
    S_A[77][25] = 4'hF;
    S_A[78][25] = 4'hF;
    S_A[79][25] = 4'hF;
    S_A[80][25] = 4'hF;
    S_A[81][25] = 4'hF;
    S_A[82][25] = 4'hF;
    S_A[83][25] = 4'hF;
    S_A[84][25] = 4'hF;
    S_A[85][25] = 4'hF;
    S_A[86][25] = 4'hF;
    S_A[87][25] = 4'hF;
    S_A[88][25] = 4'hF;
    S_A[89][25] = 4'hF;
    S_A[90][25] = 4'hF;
    S_A[91][25] = 4'hF;
    S_A[92][25] = 4'hF;
    S_A[93][25] = 4'hF;
    S_A[94][25] = 4'hF;
    S_A[95][25] = 4'hF;
    S_A[96][25] = 4'hF;
    S_A[97][25] = 4'hC;
    S_A[98][25] = 4'hC;
    S_A[99][25] = 4'hC;
    S_A[100][25] = 4'hC;
    S_A[101][25] = 4'hC;
    S_A[102][25] = 4'hC;
    S_A[103][25] = 4'hC;
    S_A[104][25] = 4'hC;
    S_A[105][25] = 4'hC;
    S_A[106][25] = 4'hC;
    S_A[107][25] = 4'hF;
    S_A[108][25] = 4'hF;
    S_A[109][25] = 4'hF;
    S_A[110][25] = 4'hF;
    S_A[111][25] = 4'hF;
    S_A[112][25] = 4'hF;
    S_A[113][25] = 4'hF;
    S_A[114][25] = 4'hF;
    S_A[0][26] = 4'hF;
    S_A[1][26] = 4'hF;
    S_A[2][26] = 4'hC;
    S_A[3][26] = 4'hC;
    S_A[4][26] = 4'hC;
    S_A[5][26] = 4'hC;
    S_A[6][26] = 4'hC;
    S_A[7][26] = 4'hC;
    S_A[8][26] = 4'hC;
    S_A[9][26] = 4'hC;
    S_A[10][26] = 4'hC;
    S_A[11][26] = 4'hC;
    S_A[12][26] = 4'hC;
    S_A[13][26] = 4'hC;
    S_A[14][26] = 4'hC;
    S_A[15][26] = 4'hC;
    S_A[16][26] = 4'hC;
    S_A[17][26] = 4'hF;
    S_A[18][26] = 4'hF;
    S_A[19][26] = 4'hF;
    S_A[20][26] = 4'hF;
    S_A[21][26] = 4'hF;
    S_A[22][26] = 4'hF;
    S_A[23][26] = 4'hF;
    S_A[24][26] = 4'hF;
    S_A[25][26] = 4'hF;
    S_A[26][26] = 4'hF;
    S_A[27][26] = 4'hF;
    S_A[28][26] = 4'hF;
    S_A[29][26] = 4'hF;
    S_A[30][26] = 4'hF;
    S_A[31][26] = 4'hF;
    S_A[32][26] = 4'hC;
    S_A[33][26] = 4'hC;
    S_A[34][26] = 4'hC;
    S_A[35][26] = 4'hC;
    S_A[36][26] = 4'hC;
    S_A[37][26] = 4'hC;
    S_A[38][26] = 4'hC;
    S_A[39][26] = 4'hC;
    S_A[40][26] = 4'hC;
    S_A[41][26] = 4'hC;
    S_A[42][26] = 4'hF;
    S_A[43][26] = 4'hF;
    S_A[44][26] = 4'hF;
    S_A[45][26] = 4'hF;
    S_A[46][26] = 4'hF;
    S_A[47][26] = 4'hF;
    S_A[48][26] = 4'hF;
    S_A[49][26] = 4'hF;
    S_A[50][26] = 4'hF;
    S_A[51][26] = 4'hF;
    S_A[52][26] = 4'hC;
    S_A[53][26] = 4'hC;
    S_A[54][26] = 4'hC;
    S_A[55][26] = 4'hC;
    S_A[56][26] = 4'hC;
    S_A[57][26] = 4'hC;
    S_A[58][26] = 4'hC;
    S_A[59][26] = 4'hC;
    S_A[60][26] = 4'hC;
    S_A[61][26] = 4'hC;
    S_A[62][26] = 4'hF;
    S_A[63][26] = 4'hF;
    S_A[64][26] = 4'hF;
    S_A[65][26] = 4'hF;
    S_A[66][26] = 4'hF;
    S_A[67][26] = 4'hF;
    S_A[68][26] = 4'hF;
    S_A[69][26] = 4'hF;
    S_A[70][26] = 4'hF;
    S_A[71][26] = 4'hF;
    S_A[72][26] = 4'hC;
    S_A[73][26] = 4'hC;
    S_A[74][26] = 4'hC;
    S_A[75][26] = 4'hC;
    S_A[76][26] = 4'hC;
    S_A[77][26] = 4'hF;
    S_A[78][26] = 4'hF;
    S_A[79][26] = 4'hF;
    S_A[80][26] = 4'hF;
    S_A[81][26] = 4'hF;
    S_A[82][26] = 4'hF;
    S_A[83][26] = 4'hF;
    S_A[84][26] = 4'hF;
    S_A[85][26] = 4'hF;
    S_A[86][26] = 4'hF;
    S_A[87][26] = 4'hF;
    S_A[88][26] = 4'hF;
    S_A[89][26] = 4'hF;
    S_A[90][26] = 4'hF;
    S_A[91][26] = 4'hF;
    S_A[92][26] = 4'hF;
    S_A[93][26] = 4'hF;
    S_A[94][26] = 4'hF;
    S_A[95][26] = 4'hF;
    S_A[96][26] = 4'hF;
    S_A[97][26] = 4'hC;
    S_A[98][26] = 4'hC;
    S_A[99][26] = 4'hC;
    S_A[100][26] = 4'hC;
    S_A[101][26] = 4'hC;
    S_A[102][26] = 4'hC;
    S_A[103][26] = 4'hC;
    S_A[104][26] = 4'hC;
    S_A[105][26] = 4'hC;
    S_A[106][26] = 4'hC;
    S_A[107][26] = 4'hF;
    S_A[108][26] = 4'hF;
    S_A[109][26] = 4'hF;
    S_A[110][26] = 4'hF;
    S_A[111][26] = 4'hF;
    S_A[112][26] = 4'hF;
    S_A[113][26] = 4'hF;
    S_A[114][26] = 4'hF;
    S_A[0][27] = 4'hF;
    S_A[1][27] = 4'hF;
    S_A[2][27] = 4'hF;
    S_A[3][27] = 4'hF;
    S_A[4][27] = 4'hF;
    S_A[5][27] = 4'hF;
    S_A[6][27] = 4'hF;
    S_A[7][27] = 4'hF;
    S_A[8][27] = 4'hF;
    S_A[9][27] = 4'hF;
    S_A[10][27] = 4'hF;
    S_A[11][27] = 4'hF;
    S_A[12][27] = 4'hF;
    S_A[13][27] = 4'hF;
    S_A[14][27] = 4'hF;
    S_A[15][27] = 4'hF;
    S_A[16][27] = 4'hF;
    S_A[17][27] = 4'hF;
    S_A[18][27] = 4'hF;
    S_A[19][27] = 4'hF;
    S_A[20][27] = 4'hF;
    S_A[21][27] = 4'hF;
    S_A[22][27] = 4'hF;
    S_A[23][27] = 4'hF;
    S_A[24][27] = 4'hF;
    S_A[25][27] = 4'hF;
    S_A[26][27] = 4'hF;
    S_A[27][27] = 4'hF;
    S_A[28][27] = 4'hF;
    S_A[29][27] = 4'hF;
    S_A[30][27] = 4'hF;
    S_A[31][27] = 4'hF;
    S_A[32][27] = 4'hF;
    S_A[33][27] = 4'hF;
    S_A[34][27] = 4'hF;
    S_A[35][27] = 4'hF;
    S_A[36][27] = 4'hF;
    S_A[37][27] = 4'hF;
    S_A[38][27] = 4'hF;
    S_A[39][27] = 4'hF;
    S_A[40][27] = 4'hF;
    S_A[41][27] = 4'hF;
    S_A[42][27] = 4'hF;
    S_A[43][27] = 4'hF;
    S_A[44][27] = 4'hF;
    S_A[45][27] = 4'hF;
    S_A[46][27] = 4'hF;
    S_A[47][27] = 4'hF;
    S_A[48][27] = 4'hF;
    S_A[49][27] = 4'hF;
    S_A[50][27] = 4'hF;
    S_A[51][27] = 4'hF;
    S_A[52][27] = 4'hF;
    S_A[53][27] = 4'hF;
    S_A[54][27] = 4'hF;
    S_A[55][27] = 4'hF;
    S_A[56][27] = 4'hF;
    S_A[57][27] = 4'hF;
    S_A[58][27] = 4'hF;
    S_A[59][27] = 4'hF;
    S_A[60][27] = 4'hF;
    S_A[61][27] = 4'hF;
    S_A[62][27] = 4'hF;
    S_A[63][27] = 4'hF;
    S_A[64][27] = 4'hF;
    S_A[65][27] = 4'hF;
    S_A[66][27] = 4'hF;
    S_A[67][27] = 4'hF;
    S_A[68][27] = 4'hF;
    S_A[69][27] = 4'hF;
    S_A[70][27] = 4'hF;
    S_A[71][27] = 4'hF;
    S_A[72][27] = 4'hF;
    S_A[73][27] = 4'hF;
    S_A[74][27] = 4'hF;
    S_A[75][27] = 4'hF;
    S_A[76][27] = 4'hF;
    S_A[77][27] = 4'hF;
    S_A[78][27] = 4'hF;
    S_A[79][27] = 4'hF;
    S_A[80][27] = 4'hF;
    S_A[81][27] = 4'hF;
    S_A[82][27] = 4'hF;
    S_A[83][27] = 4'hF;
    S_A[84][27] = 4'hF;
    S_A[85][27] = 4'hF;
    S_A[86][27] = 4'hF;
    S_A[87][27] = 4'hF;
    S_A[88][27] = 4'hF;
    S_A[89][27] = 4'hF;
    S_A[90][27] = 4'hF;
    S_A[91][27] = 4'hF;
    S_A[92][27] = 4'hF;
    S_A[93][27] = 4'hF;
    S_A[94][27] = 4'hF;
    S_A[95][27] = 4'hF;
    S_A[96][27] = 4'hF;
    S_A[97][27] = 4'hF;
    S_A[98][27] = 4'hF;
    S_A[99][27] = 4'hF;
    S_A[100][27] = 4'hF;
    S_A[101][27] = 4'hF;
    S_A[102][27] = 4'hF;
    S_A[103][27] = 4'hF;
    S_A[104][27] = 4'hF;
    S_A[105][27] = 4'hF;
    S_A[106][27] = 4'hF;
    S_A[107][27] = 4'hF;
    S_A[108][27] = 4'hF;
    S_A[109][27] = 4'hF;
    S_A[110][27] = 4'hF;
    S_A[111][27] = 4'hF;
    S_A[112][27] = 4'hF;
    S_A[113][27] = 4'hF;
    S_A[114][27] = 4'hF;
    S_A[0][28] = 4'hF;
    S_A[1][28] = 4'hF;
    S_A[2][28] = 4'hF;
    S_A[3][28] = 4'hF;
    S_A[4][28] = 4'hF;
    S_A[5][28] = 4'hF;
    S_A[6][28] = 4'hF;
    S_A[7][28] = 4'hF;
    S_A[8][28] = 4'hF;
    S_A[9][28] = 4'hF;
    S_A[10][28] = 4'hF;
    S_A[11][28] = 4'hF;
    S_A[12][28] = 4'hF;
    S_A[13][28] = 4'hF;
    S_A[14][28] = 4'hF;
    S_A[15][28] = 4'hF;
    S_A[16][28] = 4'hF;
    S_A[17][28] = 4'hF;
    S_A[18][28] = 4'hF;
    S_A[19][28] = 4'hF;
    S_A[20][28] = 4'hF;
    S_A[21][28] = 4'hF;
    S_A[22][28] = 4'hF;
    S_A[23][28] = 4'hF;
    S_A[24][28] = 4'hF;
    S_A[25][28] = 4'hF;
    S_A[26][28] = 4'hF;
    S_A[27][28] = 4'hF;
    S_A[28][28] = 4'hF;
    S_A[29][28] = 4'hF;
    S_A[30][28] = 4'hF;
    S_A[31][28] = 4'hF;
    S_A[32][28] = 4'hF;
    S_A[33][28] = 4'hF;
    S_A[34][28] = 4'hF;
    S_A[35][28] = 4'hF;
    S_A[36][28] = 4'hF;
    S_A[37][28] = 4'hF;
    S_A[38][28] = 4'hF;
    S_A[39][28] = 4'hF;
    S_A[40][28] = 4'hF;
    S_A[41][28] = 4'hF;
    S_A[42][28] = 4'hF;
    S_A[43][28] = 4'hF;
    S_A[44][28] = 4'hF;
    S_A[45][28] = 4'hF;
    S_A[46][28] = 4'hF;
    S_A[47][28] = 4'hF;
    S_A[48][28] = 4'hF;
    S_A[49][28] = 4'hF;
    S_A[50][28] = 4'hF;
    S_A[51][28] = 4'hF;
    S_A[52][28] = 4'hF;
    S_A[53][28] = 4'hF;
    S_A[54][28] = 4'hF;
    S_A[55][28] = 4'hF;
    S_A[56][28] = 4'hF;
    S_A[57][28] = 4'hF;
    S_A[58][28] = 4'hF;
    S_A[59][28] = 4'hF;
    S_A[60][28] = 4'hF;
    S_A[61][28] = 4'hF;
    S_A[62][28] = 4'hF;
    S_A[63][28] = 4'hF;
    S_A[64][28] = 4'hF;
    S_A[65][28] = 4'hF;
    S_A[66][28] = 4'hF;
    S_A[67][28] = 4'hF;
    S_A[68][28] = 4'hF;
    S_A[69][28] = 4'hF;
    S_A[70][28] = 4'hF;
    S_A[71][28] = 4'hF;
    S_A[72][28] = 4'hF;
    S_A[73][28] = 4'hF;
    S_A[74][28] = 4'hF;
    S_A[75][28] = 4'hF;
    S_A[76][28] = 4'hF;
    S_A[77][28] = 4'hF;
    S_A[78][28] = 4'hF;
    S_A[79][28] = 4'hF;
    S_A[80][28] = 4'hF;
    S_A[81][28] = 4'hF;
    S_A[82][28] = 4'hF;
    S_A[83][28] = 4'hF;
    S_A[84][28] = 4'hF;
    S_A[85][28] = 4'hF;
    S_A[86][28] = 4'hF;
    S_A[87][28] = 4'hF;
    S_A[88][28] = 4'hF;
    S_A[89][28] = 4'hF;
    S_A[90][28] = 4'hF;
    S_A[91][28] = 4'hF;
    S_A[92][28] = 4'hF;
    S_A[93][28] = 4'hF;
    S_A[94][28] = 4'hF;
    S_A[95][28] = 4'hF;
    S_A[96][28] = 4'hF;
    S_A[97][28] = 4'hF;
    S_A[98][28] = 4'hF;
    S_A[99][28] = 4'hF;
    S_A[100][28] = 4'hF;
    S_A[101][28] = 4'hF;
    S_A[102][28] = 4'hF;
    S_A[103][28] = 4'hF;
    S_A[104][28] = 4'hF;
    S_A[105][28] = 4'hF;
    S_A[106][28] = 4'hF;
    S_A[107][28] = 4'hF;
    S_A[108][28] = 4'hF;
    S_A[109][28] = 4'hF;
    S_A[110][28] = 4'hF;
    S_A[111][28] = 4'hF;
    S_A[112][28] = 4'hF;
    S_A[113][28] = 4'hF;
    S_A[114][28] = 4'hF;

// Weapon article
    W_A[0][0] = 4'hF;
    W_A[1][0] = 4'hF;
    W_A[2][0] = 4'hF;
    W_A[3][0] = 4'hF;
    W_A[4][0] = 4'hF;
    W_A[5][0] = 4'hF;
    W_A[6][0] = 4'hF;
    W_A[7][0] = 4'hF;
    W_A[8][0] = 4'hF;
    W_A[9][0] = 4'hF;
    W_A[10][0] = 4'hF;
    W_A[11][0] = 4'hF;
    W_A[12][0] = 4'hF;
    W_A[13][0] = 4'hF;
    W_A[14][0] = 4'hF;
    W_A[15][0] = 4'hF;
    W_A[16][0] = 4'hF;
    W_A[17][0] = 4'hF;
    W_A[18][0] = 4'hF;
    W_A[19][0] = 4'hF;
    W_A[20][0] = 4'hF;
    W_A[21][0] = 4'hF;
    W_A[22][0] = 4'hF;
    W_A[23][0] = 4'hF;
    W_A[24][0] = 4'hF;
    W_A[25][0] = 4'hF;
    W_A[26][0] = 4'hF;
    W_A[27][0] = 4'hF;
    W_A[28][0] = 4'hF;
    W_A[29][0] = 4'hF;
    W_A[30][0] = 4'hF;
    W_A[31][0] = 4'hF;
    W_A[32][0] = 4'hF;
    W_A[33][0] = 4'hF;
    W_A[34][0] = 4'hF;
    W_A[35][0] = 4'hF;
    W_A[36][0] = 4'hF;
    W_A[37][0] = 4'hF;
    W_A[38][0] = 4'hF;
    W_A[39][0] = 4'hF;
    W_A[40][0] = 4'hF;
    W_A[41][0] = 4'hF;
    W_A[42][0] = 4'hF;
    W_A[43][0] = 4'hF;
    W_A[44][0] = 4'hF;
    W_A[45][0] = 4'hF;
    W_A[46][0] = 4'hF;
    W_A[47][0] = 4'hF;
    W_A[48][0] = 4'hF;
    W_A[49][0] = 4'hF;
    W_A[50][0] = 4'hF;
    W_A[51][0] = 4'hF;
    W_A[52][0] = 4'hF;
    W_A[53][0] = 4'hF;
    W_A[54][0] = 4'hF;
    W_A[55][0] = 4'hF;
    W_A[56][0] = 4'hF;
    W_A[57][0] = 4'hF;
    W_A[58][0] = 4'hF;
    W_A[59][0] = 4'hF;
    W_A[60][0] = 4'hF;
    W_A[61][0] = 4'hF;
    W_A[62][0] = 4'hF;
    W_A[63][0] = 4'hF;
    W_A[64][0] = 4'hF;
    W_A[65][0] = 4'hF;
    W_A[66][0] = 4'hF;
    W_A[67][0] = 4'hF;
    W_A[68][0] = 4'hF;
    W_A[69][0] = 4'hF;
    W_A[70][0] = 4'hF;
    W_A[71][0] = 4'hF;
    W_A[72][0] = 4'hF;
    W_A[73][0] = 4'hF;
    W_A[74][0] = 4'hF;
    W_A[75][0] = 4'hF;
    W_A[76][0] = 4'hF;
    W_A[77][0] = 4'hF;
    W_A[78][0] = 4'hF;
    W_A[79][0] = 4'hF;
    W_A[80][0] = 4'hF;
    W_A[81][0] = 4'hF;
    W_A[82][0] = 4'hF;
    W_A[83][0] = 4'hF;
    W_A[84][0] = 4'hF;
    W_A[85][0] = 4'hF;
    W_A[86][0] = 4'hF;
    W_A[87][0] = 4'hF;
    W_A[88][0] = 4'hF;
    W_A[89][0] = 4'hF;
    W_A[90][0] = 4'hF;
    W_A[91][0] = 4'hF;
    W_A[92][0] = 4'hF;
    W_A[93][0] = 4'hF;
    W_A[94][0] = 4'hF;
    W_A[95][0] = 4'hF;
    W_A[96][0] = 4'hF;
    W_A[97][0] = 4'hF;
    W_A[98][0] = 4'hF;
    W_A[99][0] = 4'hF;
    W_A[100][0] = 4'hF;
    W_A[101][0] = 4'hF;
    W_A[102][0] = 4'hF;
    W_A[103][0] = 4'hF;
    W_A[104][0] = 4'hF;
    W_A[105][0] = 4'hF;
    W_A[106][0] = 4'hF;
    W_A[107][0] = 4'hF;
    W_A[0][1] = 4'hF;
    W_A[1][1] = 4'hF;
    W_A[2][1] = 4'hF;
    W_A[3][1] = 4'hF;
    W_A[4][1] = 4'hF;
    W_A[5][1] = 4'hF;
    W_A[6][1] = 4'hF;
    W_A[7][1] = 4'hF;
    W_A[8][1] = 4'hF;
    W_A[9][1] = 4'hF;
    W_A[10][1] = 4'hF;
    W_A[11][1] = 4'hF;
    W_A[12][1] = 4'hF;
    W_A[13][1] = 4'hF;
    W_A[14][1] = 4'hF;
    W_A[15][1] = 4'hF;
    W_A[16][1] = 4'hF;
    W_A[17][1] = 4'hF;
    W_A[18][1] = 4'hF;
    W_A[19][1] = 4'hF;
    W_A[20][1] = 4'hF;
    W_A[21][1] = 4'hF;
    W_A[22][1] = 4'hF;
    W_A[23][1] = 4'hF;
    W_A[24][1] = 4'hF;
    W_A[25][1] = 4'hF;
    W_A[26][1] = 4'hF;
    W_A[27][1] = 4'hF;
    W_A[28][1] = 4'hF;
    W_A[29][1] = 4'hF;
    W_A[30][1] = 4'hF;
    W_A[31][1] = 4'hF;
    W_A[32][1] = 4'hF;
    W_A[33][1] = 4'hF;
    W_A[34][1] = 4'hF;
    W_A[35][1] = 4'hF;
    W_A[36][1] = 4'hF;
    W_A[37][1] = 4'hF;
    W_A[38][1] = 4'hF;
    W_A[39][1] = 4'hF;
    W_A[40][1] = 4'hF;
    W_A[41][1] = 4'hF;
    W_A[42][1] = 4'hF;
    W_A[43][1] = 4'hF;
    W_A[44][1] = 4'hF;
    W_A[45][1] = 4'hF;
    W_A[46][1] = 4'hF;
    W_A[47][1] = 4'hF;
    W_A[48][1] = 4'hF;
    W_A[49][1] = 4'hF;
    W_A[50][1] = 4'hF;
    W_A[51][1] = 4'hF;
    W_A[52][1] = 4'hF;
    W_A[53][1] = 4'hF;
    W_A[54][1] = 4'hF;
    W_A[55][1] = 4'hF;
    W_A[56][1] = 4'hF;
    W_A[57][1] = 4'hF;
    W_A[58][1] = 4'hF;
    W_A[59][1] = 4'hF;
    W_A[60][1] = 4'hF;
    W_A[61][1] = 4'hF;
    W_A[62][1] = 4'hF;
    W_A[63][1] = 4'hF;
    W_A[64][1] = 4'hF;
    W_A[65][1] = 4'hF;
    W_A[66][1] = 4'hF;
    W_A[67][1] = 4'hF;
    W_A[68][1] = 4'hF;
    W_A[69][1] = 4'hF;
    W_A[70][1] = 4'hF;
    W_A[71][1] = 4'hF;
    W_A[72][1] = 4'hF;
    W_A[73][1] = 4'hF;
    W_A[74][1] = 4'hF;
    W_A[75][1] = 4'hF;
    W_A[76][1] = 4'hF;
    W_A[77][1] = 4'hF;
    W_A[78][1] = 4'hF;
    W_A[79][1] = 4'hF;
    W_A[80][1] = 4'hF;
    W_A[81][1] = 4'hF;
    W_A[82][1] = 4'hF;
    W_A[83][1] = 4'hF;
    W_A[84][1] = 4'hF;
    W_A[85][1] = 4'hF;
    W_A[86][1] = 4'hF;
    W_A[87][1] = 4'hF;
    W_A[88][1] = 4'hF;
    W_A[89][1] = 4'hF;
    W_A[90][1] = 4'hF;
    W_A[91][1] = 4'hF;
    W_A[92][1] = 4'hF;
    W_A[93][1] = 4'hF;
    W_A[94][1] = 4'hF;
    W_A[95][1] = 4'hF;
    W_A[96][1] = 4'hF;
    W_A[97][1] = 4'hF;
    W_A[98][1] = 4'hF;
    W_A[99][1] = 4'hF;
    W_A[100][1] = 4'hF;
    W_A[101][1] = 4'hF;
    W_A[102][1] = 4'hF;
    W_A[103][1] = 4'hF;
    W_A[104][1] = 4'hF;
    W_A[105][1] = 4'hF;
    W_A[106][1] = 4'hF;
    W_A[107][1] = 4'hF;
    W_A[0][2] = 4'hF;
    W_A[1][2] = 4'hF;
    W_A[2][2] = 4'hD;
    W_A[3][2] = 4'hC;
    W_A[4][2] = 4'hC;
    W_A[5][2] = 4'hC;
    W_A[6][2] = 4'hF;
    W_A[7][2] = 4'hF;
    W_A[8][2] = 4'hF;
    W_A[9][2] = 4'hF;
    W_A[10][2] = 4'hF;
    W_A[11][2] = 4'hF;
    W_A[12][2] = 4'hF;
    W_A[13][2] = 4'hF;
    W_A[14][2] = 4'hF;
    W_A[15][2] = 4'hF;
    W_A[16][2] = 4'hD;
    W_A[17][2] = 4'hC;
    W_A[18][2] = 4'hC;
    W_A[19][2] = 4'hC;
    W_A[20][2] = 4'hF;
    W_A[21][2] = 4'hF;
    W_A[22][2] = 4'hF;
    W_A[23][2] = 4'hF;
    W_A[24][2] = 4'hF;
    W_A[25][2] = 4'hF;
    W_A[26][2] = 4'hF;
    W_A[27][2] = 4'hF;
    W_A[28][2] = 4'hF;
    W_A[29][2] = 4'hF;
    W_A[30][2] = 4'hF;
    W_A[31][2] = 4'hF;
    W_A[32][2] = 4'hF;
    W_A[33][2] = 4'hF;
    W_A[34][2] = 4'hF;
    W_A[35][2] = 4'hF;
    W_A[36][2] = 4'hF;
    W_A[37][2] = 4'hF;
    W_A[38][2] = 4'hF;
    W_A[39][2] = 4'hF;
    W_A[40][2] = 4'hF;
    W_A[41][2] = 4'hF;
    W_A[42][2] = 4'hF;
    W_A[43][2] = 4'hF;
    W_A[44][2] = 4'hF;
    W_A[45][2] = 4'hF;
    W_A[46][2] = 4'hF;
    W_A[47][2] = 4'hF;
    W_A[48][2] = 4'hF;
    W_A[49][2] = 4'hF;
    W_A[50][2] = 4'hF;
    W_A[51][2] = 4'hF;
    W_A[52][2] = 4'hF;
    W_A[53][2] = 4'hF;
    W_A[54][2] = 4'hF;
    W_A[55][2] = 4'hF;
    W_A[56][2] = 4'hF;
    W_A[57][2] = 4'hF;
    W_A[58][2] = 4'hF;
    W_A[59][2] = 4'hF;
    W_A[60][2] = 4'hF;
    W_A[61][2] = 4'hF;
    W_A[62][2] = 4'hF;
    W_A[63][2] = 4'hF;
    W_A[64][2] = 4'hF;
    W_A[65][2] = 4'hF;
    W_A[66][2] = 4'hF;
    W_A[67][2] = 4'hF;
    W_A[68][2] = 4'hF;
    W_A[69][2] = 4'hF;
    W_A[70][2] = 4'hF;
    W_A[71][2] = 4'hF;
    W_A[72][2] = 4'hF;
    W_A[73][2] = 4'hF;
    W_A[74][2] = 4'hF;
    W_A[75][2] = 4'hF;
    W_A[76][2] = 4'hF;
    W_A[77][2] = 4'hF;
    W_A[78][2] = 4'hF;
    W_A[79][2] = 4'hF;
    W_A[80][2] = 4'hF;
    W_A[81][2] = 4'hF;
    W_A[82][2] = 4'hF;
    W_A[83][2] = 4'hF;
    W_A[84][2] = 4'hF;
    W_A[85][2] = 4'hF;
    W_A[86][2] = 4'hF;
    W_A[87][2] = 4'hF;
    W_A[88][2] = 4'hF;
    W_A[89][2] = 4'hF;
    W_A[90][2] = 4'hF;
    W_A[91][2] = 4'hF;
    W_A[92][2] = 4'hF;
    W_A[93][2] = 4'hF;
    W_A[94][2] = 4'hF;
    W_A[95][2] = 4'hF;
    W_A[96][2] = 4'hF;
    W_A[97][2] = 4'hF;
    W_A[98][2] = 4'hF;
    W_A[99][2] = 4'hF;
    W_A[100][2] = 4'hF;
    W_A[101][2] = 4'hF;
    W_A[102][2] = 4'hF;
    W_A[103][2] = 4'hF;
    W_A[104][2] = 4'hF;
    W_A[105][2] = 4'hF;
    W_A[106][2] = 4'hF;
    W_A[107][2] = 4'hF;
    W_A[0][3] = 4'hF;
    W_A[1][3] = 4'hF;
    W_A[2][3] = 4'hD;
    W_A[3][3] = 4'hC;
    W_A[4][3] = 4'hC;
    W_A[5][3] = 4'hC;
    W_A[6][3] = 4'hF;
    W_A[7][3] = 4'hF;
    W_A[8][3] = 4'hF;
    W_A[9][3] = 4'hF;
    W_A[10][3] = 4'hF;
    W_A[11][3] = 4'hF;
    W_A[12][3] = 4'hF;
    W_A[13][3] = 4'hF;
    W_A[14][3] = 4'hF;
    W_A[15][3] = 4'hF;
    W_A[16][3] = 4'hD;
    W_A[17][3] = 4'hC;
    W_A[18][3] = 4'hC;
    W_A[19][3] = 4'hC;
    W_A[20][3] = 4'hF;
    W_A[21][3] = 4'hF;
    W_A[22][3] = 4'hF;
    W_A[23][3] = 4'hF;
    W_A[24][3] = 4'hF;
    W_A[25][3] = 4'hF;
    W_A[26][3] = 4'hF;
    W_A[27][3] = 4'hF;
    W_A[28][3] = 4'hF;
    W_A[29][3] = 4'hF;
    W_A[30][3] = 4'hF;
    W_A[31][3] = 4'hF;
    W_A[32][3] = 4'hF;
    W_A[33][3] = 4'hF;
    W_A[34][3] = 4'hF;
    W_A[35][3] = 4'hF;
    W_A[36][3] = 4'hF;
    W_A[37][3] = 4'hF;
    W_A[38][3] = 4'hF;
    W_A[39][3] = 4'hF;
    W_A[40][3] = 4'hF;
    W_A[41][3] = 4'hF;
    W_A[42][3] = 4'hF;
    W_A[43][3] = 4'hF;
    W_A[44][3] = 4'hF;
    W_A[45][3] = 4'hF;
    W_A[46][3] = 4'hF;
    W_A[47][3] = 4'hF;
    W_A[48][3] = 4'hF;
    W_A[49][3] = 4'hF;
    W_A[50][3] = 4'hF;
    W_A[51][3] = 4'hF;
    W_A[52][3] = 4'hF;
    W_A[53][3] = 4'hF;
    W_A[54][3] = 4'hF;
    W_A[55][3] = 4'hF;
    W_A[56][3] = 4'hF;
    W_A[57][3] = 4'hF;
    W_A[58][3] = 4'hF;
    W_A[59][3] = 4'hF;
    W_A[60][3] = 4'hF;
    W_A[61][3] = 4'hF;
    W_A[62][3] = 4'hF;
    W_A[63][3] = 4'hF;
    W_A[64][3] = 4'hF;
    W_A[65][3] = 4'hF;
    W_A[66][3] = 4'hF;
    W_A[67][3] = 4'hF;
    W_A[68][3] = 4'hF;
    W_A[69][3] = 4'hF;
    W_A[70][3] = 4'hF;
    W_A[71][3] = 4'hF;
    W_A[72][3] = 4'hF;
    W_A[73][3] = 4'hF;
    W_A[74][3] = 4'hF;
    W_A[75][3] = 4'hF;
    W_A[76][3] = 4'hF;
    W_A[77][3] = 4'hF;
    W_A[78][3] = 4'hF;
    W_A[79][3] = 4'hF;
    W_A[80][3] = 4'hF;
    W_A[81][3] = 4'hF;
    W_A[82][3] = 4'hF;
    W_A[83][3] = 4'hF;
    W_A[84][3] = 4'hF;
    W_A[85][3] = 4'hF;
    W_A[86][3] = 4'hF;
    W_A[87][3] = 4'hF;
    W_A[88][3] = 4'hF;
    W_A[89][3] = 4'hF;
    W_A[90][3] = 4'hF;
    W_A[91][3] = 4'hF;
    W_A[92][3] = 4'hF;
    W_A[93][3] = 4'hF;
    W_A[94][3] = 4'hF;
    W_A[95][3] = 4'hF;
    W_A[96][3] = 4'hF;
    W_A[97][3] = 4'hF;
    W_A[98][3] = 4'hF;
    W_A[99][3] = 4'hF;
    W_A[100][3] = 4'hF;
    W_A[101][3] = 4'hF;
    W_A[102][3] = 4'hF;
    W_A[103][3] = 4'hF;
    W_A[104][3] = 4'hF;
    W_A[105][3] = 4'hF;
    W_A[106][3] = 4'hF;
    W_A[107][3] = 4'hF;
    W_A[0][4] = 4'hF;
    W_A[1][4] = 4'hF;
    W_A[2][4] = 4'hD;
    W_A[3][4] = 4'hC;
    W_A[4][4] = 4'hC;
    W_A[5][4] = 4'hC;
    W_A[6][4] = 4'hF;
    W_A[7][4] = 4'hF;
    W_A[8][4] = 4'hF;
    W_A[9][4] = 4'hF;
    W_A[10][4] = 4'hF;
    W_A[11][4] = 4'hF;
    W_A[12][4] = 4'hF;
    W_A[13][4] = 4'hF;
    W_A[14][4] = 4'hF;
    W_A[15][4] = 4'hF;
    W_A[16][4] = 4'hD;
    W_A[17][4] = 4'hC;
    W_A[18][4] = 4'hC;
    W_A[19][4] = 4'hC;
    W_A[20][4] = 4'hF;
    W_A[21][4] = 4'hF;
    W_A[22][4] = 4'hF;
    W_A[23][4] = 4'hF;
    W_A[24][4] = 4'hF;
    W_A[25][4] = 4'hF;
    W_A[26][4] = 4'hF;
    W_A[27][4] = 4'hF;
    W_A[28][4] = 4'hF;
    W_A[29][4] = 4'hF;
    W_A[30][4] = 4'hF;
    W_A[31][4] = 4'hF;
    W_A[32][4] = 4'hF;
    W_A[33][4] = 4'hF;
    W_A[34][4] = 4'hF;
    W_A[35][4] = 4'hF;
    W_A[36][4] = 4'hF;
    W_A[37][4] = 4'hF;
    W_A[38][4] = 4'hF;
    W_A[39][4] = 4'hF;
    W_A[40][4] = 4'hF;
    W_A[41][4] = 4'hF;
    W_A[42][4] = 4'hF;
    W_A[43][4] = 4'hF;
    W_A[44][4] = 4'hF;
    W_A[45][4] = 4'hF;
    W_A[46][4] = 4'hF;
    W_A[47][4] = 4'hF;
    W_A[48][4] = 4'hF;
    W_A[49][4] = 4'hF;
    W_A[50][4] = 4'hF;
    W_A[51][4] = 4'hF;
    W_A[52][4] = 4'hF;
    W_A[53][4] = 4'hF;
    W_A[54][4] = 4'hF;
    W_A[55][4] = 4'hF;
    W_A[56][4] = 4'hF;
    W_A[57][4] = 4'hF;
    W_A[58][4] = 4'hF;
    W_A[59][4] = 4'hF;
    W_A[60][4] = 4'hF;
    W_A[61][4] = 4'hF;
    W_A[62][4] = 4'hF;
    W_A[63][4] = 4'hF;
    W_A[64][4] = 4'hF;
    W_A[65][4] = 4'hF;
    W_A[66][4] = 4'hF;
    W_A[67][4] = 4'hF;
    W_A[68][4] = 4'hF;
    W_A[69][4] = 4'hF;
    W_A[70][4] = 4'hF;
    W_A[71][4] = 4'hF;
    W_A[72][4] = 4'hF;
    W_A[73][4] = 4'hF;
    W_A[74][4] = 4'hF;
    W_A[75][4] = 4'hF;
    W_A[76][4] = 4'hF;
    W_A[77][4] = 4'hF;
    W_A[78][4] = 4'hF;
    W_A[79][4] = 4'hF;
    W_A[80][4] = 4'hF;
    W_A[81][4] = 4'hF;
    W_A[82][4] = 4'hF;
    W_A[83][4] = 4'hF;
    W_A[84][4] = 4'hF;
    W_A[85][4] = 4'hF;
    W_A[86][4] = 4'hF;
    W_A[87][4] = 4'hF;
    W_A[88][4] = 4'hF;
    W_A[89][4] = 4'hF;
    W_A[90][4] = 4'hF;
    W_A[91][4] = 4'hF;
    W_A[92][4] = 4'hF;
    W_A[93][4] = 4'hF;
    W_A[94][4] = 4'hF;
    W_A[95][4] = 4'hF;
    W_A[96][4] = 4'hF;
    W_A[97][4] = 4'hF;
    W_A[98][4] = 4'hF;
    W_A[99][4] = 4'hF;
    W_A[100][4] = 4'hF;
    W_A[101][4] = 4'hF;
    W_A[102][4] = 4'hF;
    W_A[103][4] = 4'hF;
    W_A[104][4] = 4'hF;
    W_A[105][4] = 4'hF;
    W_A[106][4] = 4'hF;
    W_A[107][4] = 4'hF;
    W_A[0][5] = 4'hF;
    W_A[1][5] = 4'hF;
    W_A[2][5] = 4'hD;
    W_A[3][5] = 4'hC;
    W_A[4][5] = 4'hC;
    W_A[5][5] = 4'hC;
    W_A[6][5] = 4'hF;
    W_A[7][5] = 4'hF;
    W_A[8][5] = 4'hF;
    W_A[9][5] = 4'hF;
    W_A[10][5] = 4'hF;
    W_A[11][5] = 4'hF;
    W_A[12][5] = 4'hF;
    W_A[13][5] = 4'hF;
    W_A[14][5] = 4'hF;
    W_A[15][5] = 4'hF;
    W_A[16][5] = 4'hD;
    W_A[17][5] = 4'hC;
    W_A[18][5] = 4'hC;
    W_A[19][5] = 4'hC;
    W_A[20][5] = 4'hF;
    W_A[21][5] = 4'hF;
    W_A[22][5] = 4'hF;
    W_A[23][5] = 4'hF;
    W_A[24][5] = 4'hF;
    W_A[25][5] = 4'hF;
    W_A[26][5] = 4'hF;
    W_A[27][5] = 4'hF;
    W_A[28][5] = 4'hF;
    W_A[29][5] = 4'hF;
    W_A[30][5] = 4'hF;
    W_A[31][5] = 4'hF;
    W_A[32][5] = 4'hF;
    W_A[33][5] = 4'hF;
    W_A[34][5] = 4'hF;
    W_A[35][5] = 4'hF;
    W_A[36][5] = 4'hF;
    W_A[37][5] = 4'hF;
    W_A[38][5] = 4'hF;
    W_A[39][5] = 4'hF;
    W_A[40][5] = 4'hF;
    W_A[41][5] = 4'hF;
    W_A[42][5] = 4'hF;
    W_A[43][5] = 4'hF;
    W_A[44][5] = 4'hF;
    W_A[45][5] = 4'hF;
    W_A[46][5] = 4'hF;
    W_A[47][5] = 4'hF;
    W_A[48][5] = 4'hF;
    W_A[49][5] = 4'hF;
    W_A[50][5] = 4'hF;
    W_A[51][5] = 4'hF;
    W_A[52][5] = 4'hF;
    W_A[53][5] = 4'hF;
    W_A[54][5] = 4'hF;
    W_A[55][5] = 4'hF;
    W_A[56][5] = 4'hF;
    W_A[57][5] = 4'hF;
    W_A[58][5] = 4'hF;
    W_A[59][5] = 4'hF;
    W_A[60][5] = 4'hF;
    W_A[61][5] = 4'hF;
    W_A[62][5] = 4'hF;
    W_A[63][5] = 4'hF;
    W_A[64][5] = 4'hF;
    W_A[65][5] = 4'hF;
    W_A[66][5] = 4'hF;
    W_A[67][5] = 4'hF;
    W_A[68][5] = 4'hF;
    W_A[69][5] = 4'hF;
    W_A[70][5] = 4'hF;
    W_A[71][5] = 4'hF;
    W_A[72][5] = 4'hF;
    W_A[73][5] = 4'hF;
    W_A[74][5] = 4'hF;
    W_A[75][5] = 4'hF;
    W_A[76][5] = 4'hF;
    W_A[77][5] = 4'hF;
    W_A[78][5] = 4'hF;
    W_A[79][5] = 4'hF;
    W_A[80][5] = 4'hF;
    W_A[81][5] = 4'hF;
    W_A[82][5] = 4'hF;
    W_A[83][5] = 4'hF;
    W_A[84][5] = 4'hF;
    W_A[85][5] = 4'hF;
    W_A[86][5] = 4'hF;
    W_A[87][5] = 4'hF;
    W_A[88][5] = 4'hF;
    W_A[89][5] = 4'hF;
    W_A[90][5] = 4'hF;
    W_A[91][5] = 4'hF;
    W_A[92][5] = 4'hF;
    W_A[93][5] = 4'hF;
    W_A[94][5] = 4'hF;
    W_A[95][5] = 4'hF;
    W_A[96][5] = 4'hF;
    W_A[97][5] = 4'hF;
    W_A[98][5] = 4'hF;
    W_A[99][5] = 4'hF;
    W_A[100][5] = 4'hF;
    W_A[101][5] = 4'hF;
    W_A[102][5] = 4'hF;
    W_A[103][5] = 4'hF;
    W_A[104][5] = 4'hF;
    W_A[105][5] = 4'hF;
    W_A[106][5] = 4'hF;
    W_A[107][5] = 4'hF;
    W_A[0][6] = 4'hF;
    W_A[1][6] = 4'hF;
    W_A[2][6] = 4'hD;
    W_A[3][6] = 4'hC;
    W_A[4][6] = 4'hC;
    W_A[5][6] = 4'hC;
    W_A[6][6] = 4'hF;
    W_A[7][6] = 4'hF;
    W_A[8][6] = 4'hF;
    W_A[9][6] = 4'hF;
    W_A[10][6] = 4'hF;
    W_A[11][6] = 4'hF;
    W_A[12][6] = 4'hF;
    W_A[13][6] = 4'hF;
    W_A[14][6] = 4'hF;
    W_A[15][6] = 4'hF;
    W_A[16][6] = 4'hD;
    W_A[17][6] = 4'hC;
    W_A[18][6] = 4'hC;
    W_A[19][6] = 4'hC;
    W_A[20][6] = 4'hF;
    W_A[21][6] = 4'hF;
    W_A[22][6] = 4'hF;
    W_A[23][6] = 4'hF;
    W_A[24][6] = 4'hF;
    W_A[25][6] = 4'hF;
    W_A[26][6] = 4'hF;
    W_A[27][6] = 4'hC;
    W_A[28][6] = 4'hC;
    W_A[29][6] = 4'hC;
    W_A[30][6] = 4'hC;
    W_A[31][6] = 4'hC;
    W_A[32][6] = 4'hC;
    W_A[33][6] = 4'hC;
    W_A[34][6] = 4'hF;
    W_A[35][6] = 4'hF;
    W_A[36][6] = 4'hF;
    W_A[37][6] = 4'hF;
    W_A[38][6] = 4'hF;
    W_A[39][6] = 4'hF;
    W_A[40][6] = 4'hF;
    W_A[41][6] = 4'hF;
    W_A[42][6] = 4'hF;
    W_A[43][6] = 4'hF;
    W_A[44][6] = 4'hC;
    W_A[45][6] = 4'hC;
    W_A[46][6] = 4'hC;
    W_A[47][6] = 4'hC;
    W_A[48][6] = 4'hC;
    W_A[49][6] = 4'hC;
    W_A[50][6] = 4'hC;
    W_A[51][6] = 4'hC;
    W_A[52][6] = 4'hC;
    W_A[53][6] = 4'hC;
    W_A[54][6] = 4'hD;
    W_A[55][6] = 4'hF;
    W_A[56][6] = 4'hF;
    W_A[57][6] = 4'hD;
    W_A[58][6] = 4'hC;
    W_A[59][6] = 4'hC;
    W_A[60][6] = 4'hC;
    W_A[61][6] = 4'hC;
    W_A[62][6] = 4'hC;
    W_A[63][6] = 4'hC;
    W_A[64][6] = 4'hC;
    W_A[65][6] = 4'hC;
    W_A[66][6] = 4'hC;
    W_A[67][6] = 4'hC;
    W_A[68][6] = 4'hF;
    W_A[69][6] = 4'hF;
    W_A[70][6] = 4'hF;
    W_A[71][6] = 4'hF;
    W_A[72][6] = 4'hF;
    W_A[73][6] = 4'hF;
    W_A[74][6] = 4'hF;
    W_A[75][6] = 4'hF;
    W_A[76][6] = 4'hF;
    W_A[77][6] = 4'hF;
    W_A[78][6] = 4'hC;
    W_A[79][6] = 4'hC;
    W_A[80][6] = 4'hC;
    W_A[81][6] = 4'hC;
    W_A[82][6] = 4'hC;
    W_A[83][6] = 4'hC;
    W_A[84][6] = 4'hC;
    W_A[85][6] = 4'hF;
    W_A[86][6] = 4'hF;
    W_A[87][6] = 4'hF;
    W_A[88][6] = 4'hF;
    W_A[89][6] = 4'hF;
    W_A[90][6] = 4'hF;
    W_A[91][6] = 4'hD;
    W_A[92][6] = 4'hC;
    W_A[93][6] = 4'hC;
    W_A[94][6] = 4'hC;
    W_A[95][6] = 4'hC;
    W_A[96][6] = 4'hC;
    W_A[97][6] = 4'hC;
    W_A[98][6] = 4'hC;
    W_A[99][6] = 4'hC;
    W_A[100][6] = 4'hC;
    W_A[101][6] = 4'hC;
    W_A[102][6] = 4'hF;
    W_A[103][6] = 4'hF;
    W_A[104][6] = 4'hF;
    W_A[105][6] = 4'hF;
    W_A[106][6] = 4'hF;
    W_A[107][6] = 4'hF;
    W_A[0][7] = 4'hF;
    W_A[1][7] = 4'hF;
    W_A[2][7] = 4'hD;
    W_A[3][7] = 4'hC;
    W_A[4][7] = 4'hC;
    W_A[5][7] = 4'hC;
    W_A[6][7] = 4'hF;
    W_A[7][7] = 4'hF;
    W_A[8][7] = 4'hF;
    W_A[9][7] = 4'hF;
    W_A[10][7] = 4'hF;
    W_A[11][7] = 4'hF;
    W_A[12][7] = 4'hF;
    W_A[13][7] = 4'hF;
    W_A[14][7] = 4'hF;
    W_A[15][7] = 4'hF;
    W_A[16][7] = 4'hD;
    W_A[17][7] = 4'hC;
    W_A[18][7] = 4'hC;
    W_A[19][7] = 4'hC;
    W_A[20][7] = 4'hF;
    W_A[21][7] = 4'hF;
    W_A[22][7] = 4'hF;
    W_A[23][7] = 4'hF;
    W_A[24][7] = 4'hF;
    W_A[25][7] = 4'hF;
    W_A[26][7] = 4'hF;
    W_A[27][7] = 4'hC;
    W_A[28][7] = 4'hC;
    W_A[29][7] = 4'hC;
    W_A[30][7] = 4'hC;
    W_A[31][7] = 4'hC;
    W_A[32][7] = 4'hC;
    W_A[33][7] = 4'hC;
    W_A[34][7] = 4'hF;
    W_A[35][7] = 4'hF;
    W_A[36][7] = 4'hF;
    W_A[37][7] = 4'hF;
    W_A[38][7] = 4'hF;
    W_A[39][7] = 4'hF;
    W_A[40][7] = 4'hF;
    W_A[41][7] = 4'hF;
    W_A[42][7] = 4'hF;
    W_A[43][7] = 4'hF;
    W_A[44][7] = 4'hC;
    W_A[45][7] = 4'hC;
    W_A[46][7] = 4'hC;
    W_A[47][7] = 4'hC;
    W_A[48][7] = 4'hC;
    W_A[49][7] = 4'hC;
    W_A[50][7] = 4'hC;
    W_A[51][7] = 4'hC;
    W_A[52][7] = 4'hC;
    W_A[53][7] = 4'hC;
    W_A[54][7] = 4'hD;
    W_A[55][7] = 4'hF;
    W_A[56][7] = 4'hF;
    W_A[57][7] = 4'hD;
    W_A[58][7] = 4'hC;
    W_A[59][7] = 4'hC;
    W_A[60][7] = 4'hC;
    W_A[61][7] = 4'hC;
    W_A[62][7] = 4'hC;
    W_A[63][7] = 4'hC;
    W_A[64][7] = 4'hC;
    W_A[65][7] = 4'hC;
    W_A[66][7] = 4'hC;
    W_A[67][7] = 4'hC;
    W_A[68][7] = 4'hF;
    W_A[69][7] = 4'hF;
    W_A[70][7] = 4'hF;
    W_A[71][7] = 4'hF;
    W_A[72][7] = 4'hF;
    W_A[73][7] = 4'hF;
    W_A[74][7] = 4'hF;
    W_A[75][7] = 4'hF;
    W_A[76][7] = 4'hF;
    W_A[77][7] = 4'hF;
    W_A[78][7] = 4'hC;
    W_A[79][7] = 4'hC;
    W_A[80][7] = 4'hC;
    W_A[81][7] = 4'hC;
    W_A[82][7] = 4'hC;
    W_A[83][7] = 4'hC;
    W_A[84][7] = 4'hC;
    W_A[85][7] = 4'hF;
    W_A[86][7] = 4'hF;
    W_A[87][7] = 4'hF;
    W_A[88][7] = 4'hF;
    W_A[89][7] = 4'hF;
    W_A[90][7] = 4'hF;
    W_A[91][7] = 4'hD;
    W_A[92][7] = 4'hC;
    W_A[93][7] = 4'hC;
    W_A[94][7] = 4'hC;
    W_A[95][7] = 4'hC;
    W_A[96][7] = 4'hC;
    W_A[97][7] = 4'hC;
    W_A[98][7] = 4'hC;
    W_A[99][7] = 4'hC;
    W_A[100][7] = 4'hC;
    W_A[101][7] = 4'hC;
    W_A[102][7] = 4'hF;
    W_A[103][7] = 4'hF;
    W_A[104][7] = 4'hF;
    W_A[105][7] = 4'hF;
    W_A[106][7] = 4'hF;
    W_A[107][7] = 4'hF;
    W_A[0][8] = 4'hF;
    W_A[1][8] = 4'hF;
    W_A[2][8] = 4'hD;
    W_A[3][8] = 4'hC;
    W_A[4][8] = 4'hC;
    W_A[5][8] = 4'hC;
    W_A[6][8] = 4'hF;
    W_A[7][8] = 4'hF;
    W_A[8][8] = 4'hF;
    W_A[9][8] = 4'hF;
    W_A[10][8] = 4'hF;
    W_A[11][8] = 4'hF;
    W_A[12][8] = 4'hF;
    W_A[13][8] = 4'hF;
    W_A[14][8] = 4'hF;
    W_A[15][8] = 4'hF;
    W_A[16][8] = 4'hD;
    W_A[17][8] = 4'hC;
    W_A[18][8] = 4'hC;
    W_A[19][8] = 4'hC;
    W_A[20][8] = 4'hF;
    W_A[21][8] = 4'hF;
    W_A[22][8] = 4'hF;
    W_A[23][8] = 4'hF;
    W_A[24][8] = 4'hF;
    W_A[25][8] = 4'hF;
    W_A[26][8] = 4'hF;
    W_A[27][8] = 4'hC;
    W_A[28][8] = 4'hC;
    W_A[29][8] = 4'hC;
    W_A[30][8] = 4'hC;
    W_A[31][8] = 4'hC;
    W_A[32][8] = 4'hC;
    W_A[33][8] = 4'hC;
    W_A[34][8] = 4'hF;
    W_A[35][8] = 4'hF;
    W_A[36][8] = 4'hF;
    W_A[37][8] = 4'hF;
    W_A[38][8] = 4'hF;
    W_A[39][8] = 4'hF;
    W_A[40][8] = 4'hF;
    W_A[41][8] = 4'hF;
    W_A[42][8] = 4'hF;
    W_A[43][8] = 4'hF;
    W_A[44][8] = 4'hC;
    W_A[45][8] = 4'hC;
    W_A[46][8] = 4'hC;
    W_A[47][8] = 4'hC;
    W_A[48][8] = 4'hC;
    W_A[49][8] = 4'hC;
    W_A[50][8] = 4'hC;
    W_A[51][8] = 4'hC;
    W_A[52][8] = 4'hC;
    W_A[53][8] = 4'hC;
    W_A[54][8] = 4'hD;
    W_A[55][8] = 4'hF;
    W_A[56][8] = 4'hF;
    W_A[57][8] = 4'hD;
    W_A[58][8] = 4'hC;
    W_A[59][8] = 4'hC;
    W_A[60][8] = 4'hC;
    W_A[61][8] = 4'hC;
    W_A[62][8] = 4'hC;
    W_A[63][8] = 4'hC;
    W_A[64][8] = 4'hC;
    W_A[65][8] = 4'hC;
    W_A[66][8] = 4'hC;
    W_A[67][8] = 4'hC;
    W_A[68][8] = 4'hF;
    W_A[69][8] = 4'hF;
    W_A[70][8] = 4'hF;
    W_A[71][8] = 4'hF;
    W_A[72][8] = 4'hF;
    W_A[73][8] = 4'hF;
    W_A[74][8] = 4'hF;
    W_A[75][8] = 4'hF;
    W_A[76][8] = 4'hF;
    W_A[77][8] = 4'hF;
    W_A[78][8] = 4'hC;
    W_A[79][8] = 4'hC;
    W_A[80][8] = 4'hC;
    W_A[81][8] = 4'hC;
    W_A[82][8] = 4'hC;
    W_A[83][8] = 4'hC;
    W_A[84][8] = 4'hC;
    W_A[85][8] = 4'hF;
    W_A[86][8] = 4'hF;
    W_A[87][8] = 4'hF;
    W_A[88][8] = 4'hF;
    W_A[89][8] = 4'hF;
    W_A[90][8] = 4'hF;
    W_A[91][8] = 4'hD;
    W_A[92][8] = 4'hC;
    W_A[93][8] = 4'hC;
    W_A[94][8] = 4'hC;
    W_A[95][8] = 4'hC;
    W_A[96][8] = 4'hC;
    W_A[97][8] = 4'hC;
    W_A[98][8] = 4'hC;
    W_A[99][8] = 4'hC;
    W_A[100][8] = 4'hC;
    W_A[101][8] = 4'hC;
    W_A[102][8] = 4'hF;
    W_A[103][8] = 4'hF;
    W_A[104][8] = 4'hF;
    W_A[105][8] = 4'hF;
    W_A[106][8] = 4'hF;
    W_A[107][8] = 4'hF;
    W_A[0][9] = 4'hF;
    W_A[1][9] = 4'hF;
    W_A[2][9] = 4'hD;
    W_A[3][9] = 4'hC;
    W_A[4][9] = 4'hC;
    W_A[5][9] = 4'hC;
    W_A[6][9] = 4'hF;
    W_A[7][9] = 4'hF;
    W_A[8][9] = 4'hF;
    W_A[9][9] = 4'hE;
    W_A[10][9] = 4'hD;
    W_A[11][9] = 4'hD;
    W_A[12][9] = 4'hD;
    W_A[13][9] = 4'hF;
    W_A[14][9] = 4'hF;
    W_A[15][9] = 4'hF;
    W_A[16][9] = 4'hD;
    W_A[17][9] = 4'hC;
    W_A[18][9] = 4'hC;
    W_A[19][9] = 4'hC;
    W_A[20][9] = 4'hF;
    W_A[21][9] = 4'hF;
    W_A[22][9] = 4'hF;
    W_A[23][9] = 4'hD;
    W_A[24][9] = 4'hC;
    W_A[25][9] = 4'hC;
    W_A[26][9] = 4'hC;
    W_A[27][9] = 4'hF;
    W_A[28][9] = 4'hF;
    W_A[29][9] = 4'hF;
    W_A[30][9] = 4'hD;
    W_A[31][9] = 4'hC;
    W_A[32][9] = 4'hC;
    W_A[33][9] = 4'hC;
    W_A[34][9] = 4'hC;
    W_A[35][9] = 4'hC;
    W_A[36][9] = 4'hC;
    W_A[37][9] = 4'hD;
    W_A[38][9] = 4'hF;
    W_A[39][9] = 4'hF;
    W_A[40][9] = 4'hD;
    W_A[41][9] = 4'hC;
    W_A[42][9] = 4'hC;
    W_A[43][9] = 4'hC;
    W_A[44][9] = 4'hF;
    W_A[45][9] = 4'hF;
    W_A[46][9] = 4'hF;
    W_A[47][9] = 4'hF;
    W_A[48][9] = 4'hF;
    W_A[49][9] = 4'hF;
    W_A[50][9] = 4'hF;
    W_A[51][9] = 4'hC;
    W_A[52][9] = 4'hC;
    W_A[53][9] = 4'hC;
    W_A[54][9] = 4'hD;
    W_A[55][9] = 4'hF;
    W_A[56][9] = 4'hF;
    W_A[57][9] = 4'hD;
    W_A[58][9] = 4'hC;
    W_A[59][9] = 4'hC;
    W_A[60][9] = 4'hC;
    W_A[61][9] = 4'hF;
    W_A[62][9] = 4'hF;
    W_A[63][9] = 4'hF;
    W_A[64][9] = 4'hF;
    W_A[65][9] = 4'hF;
    W_A[66][9] = 4'hF;
    W_A[67][9] = 4'hF;
    W_A[68][9] = 4'hC;
    W_A[69][9] = 4'hC;
    W_A[70][9] = 4'hC;
    W_A[71][9] = 4'hD;
    W_A[72][9] = 4'hF;
    W_A[73][9] = 4'hF;
    W_A[74][9] = 4'hD;
    W_A[75][9] = 4'hC;
    W_A[76][9] = 4'hC;
    W_A[77][9] = 4'hC;
    W_A[78][9] = 4'hF;
    W_A[79][9] = 4'hF;
    W_A[80][9] = 4'hF;
    W_A[81][9] = 4'hF;
    W_A[82][9] = 4'hF;
    W_A[83][9] = 4'hF;
    W_A[84][9] = 4'hF;
    W_A[85][9] = 4'hC;
    W_A[86][9] = 4'hC;
    W_A[87][9] = 4'hC;
    W_A[88][9] = 4'hD;
    W_A[89][9] = 4'hF;
    W_A[90][9] = 4'hF;
    W_A[91][9] = 4'hD;
    W_A[92][9] = 4'hC;
    W_A[93][9] = 4'hC;
    W_A[94][9] = 4'hC;
    W_A[95][9] = 4'hD;
    W_A[96][9] = 4'hD;
    W_A[97][9] = 4'hD;
    W_A[98][9] = 4'hD;
    W_A[99][9] = 4'hD;
    W_A[100][9] = 4'hD;
    W_A[101][9] = 4'hD;
    W_A[102][9] = 4'hD;
    W_A[103][9] = 4'hD;
    W_A[104][9] = 4'hD;
    W_A[105][9] = 4'hE;
    W_A[106][9] = 4'hF;
    W_A[107][9] = 4'hF;
    W_A[0][10] = 4'hF;
    W_A[1][10] = 4'hF;
    W_A[2][10] = 4'hD;
    W_A[3][10] = 4'hC;
    W_A[4][10] = 4'hC;
    W_A[5][10] = 4'hC;
    W_A[6][10] = 4'hF;
    W_A[7][10] = 4'hF;
    W_A[8][10] = 4'hF;
    W_A[9][10] = 4'hD;
    W_A[10][10] = 4'hC;
    W_A[11][10] = 4'hC;
    W_A[12][10] = 4'hC;
    W_A[13][10] = 4'hF;
    W_A[14][10] = 4'hF;
    W_A[15][10] = 4'hF;
    W_A[16][10] = 4'hD;
    W_A[17][10] = 4'hC;
    W_A[18][10] = 4'hC;
    W_A[19][10] = 4'hC;
    W_A[20][10] = 4'hF;
    W_A[21][10] = 4'hF;
    W_A[22][10] = 4'hF;
    W_A[23][10] = 4'hD;
    W_A[24][10] = 4'hC;
    W_A[25][10] = 4'hC;
    W_A[26][10] = 4'hC;
    W_A[27][10] = 4'hF;
    W_A[28][10] = 4'hF;
    W_A[29][10] = 4'hF;
    W_A[30][10] = 4'hD;
    W_A[31][10] = 4'hC;
    W_A[32][10] = 4'hC;
    W_A[33][10] = 4'hC;
    W_A[34][10] = 4'hC;
    W_A[35][10] = 4'hC;
    W_A[36][10] = 4'hC;
    W_A[37][10] = 4'hD;
    W_A[38][10] = 4'hF;
    W_A[39][10] = 4'hF;
    W_A[40][10] = 4'hD;
    W_A[41][10] = 4'hC;
    W_A[42][10] = 4'hC;
    W_A[43][10] = 4'hC;
    W_A[44][10] = 4'hF;
    W_A[45][10] = 4'hF;
    W_A[46][10] = 4'hF;
    W_A[47][10] = 4'hF;
    W_A[48][10] = 4'hF;
    W_A[49][10] = 4'hF;
    W_A[50][10] = 4'hF;
    W_A[51][10] = 4'hC;
    W_A[52][10] = 4'hC;
    W_A[53][10] = 4'hC;
    W_A[54][10] = 4'hD;
    W_A[55][10] = 4'hF;
    W_A[56][10] = 4'hF;
    W_A[57][10] = 4'hD;
    W_A[58][10] = 4'hC;
    W_A[59][10] = 4'hC;
    W_A[60][10] = 4'hC;
    W_A[61][10] = 4'hF;
    W_A[62][10] = 4'hF;
    W_A[63][10] = 4'hF;
    W_A[64][10] = 4'hF;
    W_A[65][10] = 4'hF;
    W_A[66][10] = 4'hF;
    W_A[67][10] = 4'hF;
    W_A[68][10] = 4'hC;
    W_A[69][10] = 4'hC;
    W_A[70][10] = 4'hC;
    W_A[71][10] = 4'hD;
    W_A[72][10] = 4'hF;
    W_A[73][10] = 4'hF;
    W_A[74][10] = 4'hD;
    W_A[75][10] = 4'hC;
    W_A[76][10] = 4'hC;
    W_A[77][10] = 4'hC;
    W_A[78][10] = 4'hF;
    W_A[79][10] = 4'hF;
    W_A[80][10] = 4'hF;
    W_A[81][10] = 4'hF;
    W_A[82][10] = 4'hF;
    W_A[83][10] = 4'hF;
    W_A[84][10] = 4'hF;
    W_A[85][10] = 4'hC;
    W_A[86][10] = 4'hC;
    W_A[87][10] = 4'hC;
    W_A[88][10] = 4'hD;
    W_A[89][10] = 4'hF;
    W_A[90][10] = 4'hF;
    W_A[91][10] = 4'hD;
    W_A[92][10] = 4'hC;
    W_A[93][10] = 4'hC;
    W_A[94][10] = 4'hC;
    W_A[95][10] = 4'hF;
    W_A[96][10] = 4'hF;
    W_A[97][10] = 4'hF;
    W_A[98][10] = 4'hF;
    W_A[99][10] = 4'hF;
    W_A[100][10] = 4'hF;
    W_A[101][10] = 4'hF;
    W_A[102][10] = 4'hC;
    W_A[103][10] = 4'hC;
    W_A[104][10] = 4'hC;
    W_A[105][10] = 4'hD;
    W_A[106][10] = 4'hF;
    W_A[107][10] = 4'hF;
    W_A[0][11] = 4'hF;
    W_A[1][11] = 4'hF;
    W_A[2][11] = 4'hD;
    W_A[3][11] = 4'hC;
    W_A[4][11] = 4'hC;
    W_A[5][11] = 4'hC;
    W_A[6][11] = 4'hF;
    W_A[7][11] = 4'hF;
    W_A[8][11] = 4'hF;
    W_A[9][11] = 4'hD;
    W_A[10][11] = 4'hC;
    W_A[11][11] = 4'hC;
    W_A[12][11] = 4'hC;
    W_A[13][11] = 4'hF;
    W_A[14][11] = 4'hF;
    W_A[15][11] = 4'hF;
    W_A[16][11] = 4'hD;
    W_A[17][11] = 4'hC;
    W_A[18][11] = 4'hC;
    W_A[19][11] = 4'hC;
    W_A[20][11] = 4'hF;
    W_A[21][11] = 4'hF;
    W_A[22][11] = 4'hF;
    W_A[23][11] = 4'hD;
    W_A[24][11] = 4'hC;
    W_A[25][11] = 4'hC;
    W_A[26][11] = 4'hC;
    W_A[27][11] = 4'hF;
    W_A[28][11] = 4'hF;
    W_A[29][11] = 4'hF;
    W_A[30][11] = 4'hD;
    W_A[31][11] = 4'hC;
    W_A[32][11] = 4'hC;
    W_A[33][11] = 4'hC;
    W_A[34][11] = 4'hC;
    W_A[35][11] = 4'hC;
    W_A[36][11] = 4'hC;
    W_A[37][11] = 4'hD;
    W_A[38][11] = 4'hF;
    W_A[39][11] = 4'hF;
    W_A[40][11] = 4'hD;
    W_A[41][11] = 4'hC;
    W_A[42][11] = 4'hC;
    W_A[43][11] = 4'hC;
    W_A[44][11] = 4'hF;
    W_A[45][11] = 4'hF;
    W_A[46][11] = 4'hF;
    W_A[47][11] = 4'hF;
    W_A[48][11] = 4'hF;
    W_A[49][11] = 4'hF;
    W_A[50][11] = 4'hF;
    W_A[51][11] = 4'hC;
    W_A[52][11] = 4'hC;
    W_A[53][11] = 4'hC;
    W_A[54][11] = 4'hD;
    W_A[55][11] = 4'hF;
    W_A[56][11] = 4'hF;
    W_A[57][11] = 4'hD;
    W_A[58][11] = 4'hC;
    W_A[59][11] = 4'hC;
    W_A[60][11] = 4'hC;
    W_A[61][11] = 4'hF;
    W_A[62][11] = 4'hF;
    W_A[63][11] = 4'hF;
    W_A[64][11] = 4'hF;
    W_A[65][11] = 4'hF;
    W_A[66][11] = 4'hF;
    W_A[67][11] = 4'hF;
    W_A[68][11] = 4'hC;
    W_A[69][11] = 4'hC;
    W_A[70][11] = 4'hC;
    W_A[71][11] = 4'hD;
    W_A[72][11] = 4'hF;
    W_A[73][11] = 4'hF;
    W_A[74][11] = 4'hD;
    W_A[75][11] = 4'hC;
    W_A[76][11] = 4'hC;
    W_A[77][11] = 4'hC;
    W_A[78][11] = 4'hF;
    W_A[79][11] = 4'hF;
    W_A[80][11] = 4'hF;
    W_A[81][11] = 4'hF;
    W_A[82][11] = 4'hF;
    W_A[83][11] = 4'hF;
    W_A[84][11] = 4'hF;
    W_A[85][11] = 4'hC;
    W_A[86][11] = 4'hC;
    W_A[87][11] = 4'hC;
    W_A[88][11] = 4'hD;
    W_A[89][11] = 4'hF;
    W_A[90][11] = 4'hF;
    W_A[91][11] = 4'hD;
    W_A[92][11] = 4'hC;
    W_A[93][11] = 4'hC;
    W_A[94][11] = 4'hC;
    W_A[95][11] = 4'hF;
    W_A[96][11] = 4'hF;
    W_A[97][11] = 4'hF;
    W_A[98][11] = 4'hF;
    W_A[99][11] = 4'hF;
    W_A[100][11] = 4'hF;
    W_A[101][11] = 4'hF;
    W_A[102][11] = 4'hC;
    W_A[103][11] = 4'hC;
    W_A[104][11] = 4'hC;
    W_A[105][11] = 4'hD;
    W_A[106][11] = 4'hF;
    W_A[107][11] = 4'hF;
    W_A[0][12] = 4'hF;
    W_A[1][12] = 4'hF;
    W_A[2][12] = 4'hD;
    W_A[3][12] = 4'hC;
    W_A[4][12] = 4'hC;
    W_A[5][12] = 4'hC;
    W_A[6][12] = 4'hF;
    W_A[7][12] = 4'hF;
    W_A[8][12] = 4'hF;
    W_A[9][12] = 4'hD;
    W_A[10][12] = 4'hC;
    W_A[11][12] = 4'hC;
    W_A[12][12] = 4'hC;
    W_A[13][12] = 4'hF;
    W_A[14][12] = 4'hF;
    W_A[15][12] = 4'hF;
    W_A[16][12] = 4'hD;
    W_A[17][12] = 4'hC;
    W_A[18][12] = 4'hC;
    W_A[19][12] = 4'hC;
    W_A[20][12] = 4'hF;
    W_A[21][12] = 4'hF;
    W_A[22][12] = 4'hF;
    W_A[23][12] = 4'hD;
    W_A[24][12] = 4'hC;
    W_A[25][12] = 4'hC;
    W_A[26][12] = 4'hC;
    W_A[27][12] = 4'hF;
    W_A[28][12] = 4'hF;
    W_A[29][12] = 4'hF;
    W_A[30][12] = 4'hD;
    W_A[31][12] = 4'hC;
    W_A[32][12] = 4'hC;
    W_A[33][12] = 4'hC;
    W_A[34][12] = 4'hC;
    W_A[35][12] = 4'hC;
    W_A[36][12] = 4'hC;
    W_A[37][12] = 4'hD;
    W_A[38][12] = 4'hF;
    W_A[39][12] = 4'hF;
    W_A[40][12] = 4'hD;
    W_A[41][12] = 4'hC;
    W_A[42][12] = 4'hC;
    W_A[43][12] = 4'hC;
    W_A[44][12] = 4'hF;
    W_A[45][12] = 4'hF;
    W_A[46][12] = 4'hF;
    W_A[47][12] = 4'hF;
    W_A[48][12] = 4'hF;
    W_A[49][12] = 4'hF;
    W_A[50][12] = 4'hF;
    W_A[51][12] = 4'hC;
    W_A[52][12] = 4'hC;
    W_A[53][12] = 4'hC;
    W_A[54][12] = 4'hD;
    W_A[55][12] = 4'hF;
    W_A[56][12] = 4'hF;
    W_A[57][12] = 4'hD;
    W_A[58][12] = 4'hC;
    W_A[59][12] = 4'hC;
    W_A[60][12] = 4'hC;
    W_A[61][12] = 4'hF;
    W_A[62][12] = 4'hF;
    W_A[63][12] = 4'hF;
    W_A[64][12] = 4'hF;
    W_A[65][12] = 4'hF;
    W_A[66][12] = 4'hF;
    W_A[67][12] = 4'hF;
    W_A[68][12] = 4'hC;
    W_A[69][12] = 4'hC;
    W_A[70][12] = 4'hC;
    W_A[71][12] = 4'hD;
    W_A[72][12] = 4'hF;
    W_A[73][12] = 4'hF;
    W_A[74][12] = 4'hD;
    W_A[75][12] = 4'hC;
    W_A[76][12] = 4'hC;
    W_A[77][12] = 4'hC;
    W_A[78][12] = 4'hF;
    W_A[79][12] = 4'hF;
    W_A[80][12] = 4'hF;
    W_A[81][12] = 4'hF;
    W_A[82][12] = 4'hF;
    W_A[83][12] = 4'hF;
    W_A[84][12] = 4'hF;
    W_A[85][12] = 4'hC;
    W_A[86][12] = 4'hC;
    W_A[87][12] = 4'hC;
    W_A[88][12] = 4'hD;
    W_A[89][12] = 4'hF;
    W_A[90][12] = 4'hF;
    W_A[91][12] = 4'hD;
    W_A[92][12] = 4'hC;
    W_A[93][12] = 4'hC;
    W_A[94][12] = 4'hC;
    W_A[95][12] = 4'hF;
    W_A[96][12] = 4'hF;
    W_A[97][12] = 4'hF;
    W_A[98][12] = 4'hF;
    W_A[99][12] = 4'hF;
    W_A[100][12] = 4'hF;
    W_A[101][12] = 4'hF;
    W_A[102][12] = 4'hC;
    W_A[103][12] = 4'hC;
    W_A[104][12] = 4'hC;
    W_A[105][12] = 4'hD;
    W_A[106][12] = 4'hF;
    W_A[107][12] = 4'hF;
    W_A[0][13] = 4'hF;
    W_A[1][13] = 4'hF;
    W_A[2][13] = 4'hD;
    W_A[3][13] = 4'hC;
    W_A[4][13] = 4'hC;
    W_A[5][13] = 4'hC;
    W_A[6][13] = 4'hF;
    W_A[7][13] = 4'hF;
    W_A[8][13] = 4'hF;
    W_A[9][13] = 4'hD;
    W_A[10][13] = 4'hC;
    W_A[11][13] = 4'hC;
    W_A[12][13] = 4'hC;
    W_A[13][13] = 4'hF;
    W_A[14][13] = 4'hF;
    W_A[15][13] = 4'hF;
    W_A[16][13] = 4'hD;
    W_A[17][13] = 4'hC;
    W_A[18][13] = 4'hC;
    W_A[19][13] = 4'hC;
    W_A[20][13] = 4'hF;
    W_A[21][13] = 4'hF;
    W_A[22][13] = 4'hF;
    W_A[23][13] = 4'hD;
    W_A[24][13] = 4'hC;
    W_A[25][13] = 4'hC;
    W_A[26][13] = 4'hC;
    W_A[27][13] = 4'hC;
    W_A[28][13] = 4'hC;
    W_A[29][13] = 4'hC;
    W_A[30][13] = 4'hD;
    W_A[31][13] = 4'hF;
    W_A[32][13] = 4'hF;
    W_A[33][13] = 4'hF;
    W_A[34][13] = 4'hF;
    W_A[35][13] = 4'hF;
    W_A[36][13] = 4'hF;
    W_A[37][13] = 4'hF;
    W_A[38][13] = 4'hF;
    W_A[39][13] = 4'hF;
    W_A[40][13] = 4'hD;
    W_A[41][13] = 4'hC;
    W_A[42][13] = 4'hC;
    W_A[43][13] = 4'hC;
    W_A[44][13] = 4'hF;
    W_A[45][13] = 4'hF;
    W_A[46][13] = 4'hF;
    W_A[47][13] = 4'hF;
    W_A[48][13] = 4'hF;
    W_A[49][13] = 4'hF;
    W_A[50][13] = 4'hF;
    W_A[51][13] = 4'hC;
    W_A[52][13] = 4'hC;
    W_A[53][13] = 4'hC;
    W_A[54][13] = 4'hD;
    W_A[55][13] = 4'hF;
    W_A[56][13] = 4'hF;
    W_A[57][13] = 4'hD;
    W_A[58][13] = 4'hC;
    W_A[59][13] = 4'hC;
    W_A[60][13] = 4'hC;
    W_A[61][13] = 4'hF;
    W_A[62][13] = 4'hF;
    W_A[63][13] = 4'hF;
    W_A[64][13] = 4'hF;
    W_A[65][13] = 4'hF;
    W_A[66][13] = 4'hF;
    W_A[67][13] = 4'hF;
    W_A[68][13] = 4'hC;
    W_A[69][13] = 4'hC;
    W_A[70][13] = 4'hC;
    W_A[71][13] = 4'hD;
    W_A[72][13] = 4'hF;
    W_A[73][13] = 4'hF;
    W_A[74][13] = 4'hD;
    W_A[75][13] = 4'hC;
    W_A[76][13] = 4'hC;
    W_A[77][13] = 4'hC;
    W_A[78][13] = 4'hF;
    W_A[79][13] = 4'hF;
    W_A[80][13] = 4'hF;
    W_A[81][13] = 4'hF;
    W_A[82][13] = 4'hF;
    W_A[83][13] = 4'hF;
    W_A[84][13] = 4'hF;
    W_A[85][13] = 4'hC;
    W_A[86][13] = 4'hC;
    W_A[87][13] = 4'hC;
    W_A[88][13] = 4'hD;
    W_A[89][13] = 4'hF;
    W_A[90][13] = 4'hF;
    W_A[91][13] = 4'hD;
    W_A[92][13] = 4'hC;
    W_A[93][13] = 4'hC;
    W_A[94][13] = 4'hC;
    W_A[95][13] = 4'hF;
    W_A[96][13] = 4'hF;
    W_A[97][13] = 4'hF;
    W_A[98][13] = 4'hF;
    W_A[99][13] = 4'hF;
    W_A[100][13] = 4'hF;
    W_A[101][13] = 4'hF;
    W_A[102][13] = 4'hC;
    W_A[103][13] = 4'hC;
    W_A[104][13] = 4'hC;
    W_A[105][13] = 4'hD;
    W_A[106][13] = 4'hF;
    W_A[107][13] = 4'hF;
    W_A[0][14] = 4'hF;
    W_A[1][14] = 4'hF;
    W_A[2][14] = 4'hD;
    W_A[3][14] = 4'hC;
    W_A[4][14] = 4'hC;
    W_A[5][14] = 4'hC;
    W_A[6][14] = 4'hF;
    W_A[7][14] = 4'hF;
    W_A[8][14] = 4'hF;
    W_A[9][14] = 4'hD;
    W_A[10][14] = 4'hC;
    W_A[11][14] = 4'hC;
    W_A[12][14] = 4'hC;
    W_A[13][14] = 4'hF;
    W_A[14][14] = 4'hF;
    W_A[15][14] = 4'hF;
    W_A[16][14] = 4'hD;
    W_A[17][14] = 4'hC;
    W_A[18][14] = 4'hC;
    W_A[19][14] = 4'hC;
    W_A[20][14] = 4'hF;
    W_A[21][14] = 4'hF;
    W_A[22][14] = 4'hF;
    W_A[23][14] = 4'hD;
    W_A[24][14] = 4'hC;
    W_A[25][14] = 4'hC;
    W_A[26][14] = 4'hC;
    W_A[27][14] = 4'hC;
    W_A[28][14] = 4'hC;
    W_A[29][14] = 4'hC;
    W_A[30][14] = 4'hD;
    W_A[31][14] = 4'hF;
    W_A[32][14] = 4'hF;
    W_A[33][14] = 4'hF;
    W_A[34][14] = 4'hF;
    W_A[35][14] = 4'hF;
    W_A[36][14] = 4'hF;
    W_A[37][14] = 4'hF;
    W_A[38][14] = 4'hF;
    W_A[39][14] = 4'hF;
    W_A[40][14] = 4'hD;
    W_A[41][14] = 4'hC;
    W_A[42][14] = 4'hC;
    W_A[43][14] = 4'hC;
    W_A[44][14] = 4'hF;
    W_A[45][14] = 4'hF;
    W_A[46][14] = 4'hF;
    W_A[47][14] = 4'hF;
    W_A[48][14] = 4'hF;
    W_A[49][14] = 4'hF;
    W_A[50][14] = 4'hF;
    W_A[51][14] = 4'hC;
    W_A[52][14] = 4'hC;
    W_A[53][14] = 4'hC;
    W_A[54][14] = 4'hD;
    W_A[55][14] = 4'hF;
    W_A[56][14] = 4'hF;
    W_A[57][14] = 4'hD;
    W_A[58][14] = 4'hC;
    W_A[59][14] = 4'hC;
    W_A[60][14] = 4'hC;
    W_A[61][14] = 4'hF;
    W_A[62][14] = 4'hF;
    W_A[63][14] = 4'hF;
    W_A[64][14] = 4'hF;
    W_A[65][14] = 4'hF;
    W_A[66][14] = 4'hF;
    W_A[67][14] = 4'hF;
    W_A[68][14] = 4'hC;
    W_A[69][14] = 4'hC;
    W_A[70][14] = 4'hC;
    W_A[71][14] = 4'hD;
    W_A[72][14] = 4'hF;
    W_A[73][14] = 4'hF;
    W_A[74][14] = 4'hD;
    W_A[75][14] = 4'hC;
    W_A[76][14] = 4'hC;
    W_A[77][14] = 4'hC;
    W_A[78][14] = 4'hF;
    W_A[79][14] = 4'hF;
    W_A[80][14] = 4'hF;
    W_A[81][14] = 4'hF;
    W_A[82][14] = 4'hF;
    W_A[83][14] = 4'hF;
    W_A[84][14] = 4'hF;
    W_A[85][14] = 4'hC;
    W_A[86][14] = 4'hC;
    W_A[87][14] = 4'hC;
    W_A[88][14] = 4'hD;
    W_A[89][14] = 4'hF;
    W_A[90][14] = 4'hF;
    W_A[91][14] = 4'hD;
    W_A[92][14] = 4'hC;
    W_A[93][14] = 4'hC;
    W_A[94][14] = 4'hC;
    W_A[95][14] = 4'hF;
    W_A[96][14] = 4'hF;
    W_A[97][14] = 4'hF;
    W_A[98][14] = 4'hF;
    W_A[99][14] = 4'hF;
    W_A[100][14] = 4'hF;
    W_A[101][14] = 4'hF;
    W_A[102][14] = 4'hC;
    W_A[103][14] = 4'hC;
    W_A[104][14] = 4'hC;
    W_A[105][14] = 4'hD;
    W_A[106][14] = 4'hF;
    W_A[107][14] = 4'hF;
    W_A[0][15] = 4'hF;
    W_A[1][15] = 4'hF;
    W_A[2][15] = 4'hD;
    W_A[3][15] = 4'hC;
    W_A[4][15] = 4'hC;
    W_A[5][15] = 4'hC;
    W_A[6][15] = 4'hF;
    W_A[7][15] = 4'hF;
    W_A[8][15] = 4'hF;
    W_A[9][15] = 4'hD;
    W_A[10][15] = 4'hC;
    W_A[11][15] = 4'hC;
    W_A[12][15] = 4'hC;
    W_A[13][15] = 4'hF;
    W_A[14][15] = 4'hF;
    W_A[15][15] = 4'hF;
    W_A[16][15] = 4'hD;
    W_A[17][15] = 4'hC;
    W_A[18][15] = 4'hC;
    W_A[19][15] = 4'hC;
    W_A[20][15] = 4'hF;
    W_A[21][15] = 4'hF;
    W_A[22][15] = 4'hF;
    W_A[23][15] = 4'hD;
    W_A[24][15] = 4'hC;
    W_A[25][15] = 4'hC;
    W_A[26][15] = 4'hC;
    W_A[27][15] = 4'hC;
    W_A[28][15] = 4'hC;
    W_A[29][15] = 4'hC;
    W_A[30][15] = 4'hD;
    W_A[31][15] = 4'hF;
    W_A[32][15] = 4'hF;
    W_A[33][15] = 4'hF;
    W_A[34][15] = 4'hF;
    W_A[35][15] = 4'hF;
    W_A[36][15] = 4'hF;
    W_A[37][15] = 4'hF;
    W_A[38][15] = 4'hF;
    W_A[39][15] = 4'hF;
    W_A[40][15] = 4'hD;
    W_A[41][15] = 4'hC;
    W_A[42][15] = 4'hC;
    W_A[43][15] = 4'hC;
    W_A[44][15] = 4'hF;
    W_A[45][15] = 4'hF;
    W_A[46][15] = 4'hF;
    W_A[47][15] = 4'hF;
    W_A[48][15] = 4'hF;
    W_A[49][15] = 4'hF;
    W_A[50][15] = 4'hF;
    W_A[51][15] = 4'hC;
    W_A[52][15] = 4'hC;
    W_A[53][15] = 4'hC;
    W_A[54][15] = 4'hD;
    W_A[55][15] = 4'hF;
    W_A[56][15] = 4'hF;
    W_A[57][15] = 4'hD;
    W_A[58][15] = 4'hC;
    W_A[59][15] = 4'hC;
    W_A[60][15] = 4'hC;
    W_A[61][15] = 4'hF;
    W_A[62][15] = 4'hF;
    W_A[63][15] = 4'hF;
    W_A[64][15] = 4'hF;
    W_A[65][15] = 4'hF;
    W_A[66][15] = 4'hF;
    W_A[67][15] = 4'hF;
    W_A[68][15] = 4'hC;
    W_A[69][15] = 4'hC;
    W_A[70][15] = 4'hC;
    W_A[71][15] = 4'hD;
    W_A[72][15] = 4'hF;
    W_A[73][15] = 4'hF;
    W_A[74][15] = 4'hD;
    W_A[75][15] = 4'hC;
    W_A[76][15] = 4'hC;
    W_A[77][15] = 4'hC;
    W_A[78][15] = 4'hF;
    W_A[79][15] = 4'hF;
    W_A[80][15] = 4'hF;
    W_A[81][15] = 4'hF;
    W_A[82][15] = 4'hF;
    W_A[83][15] = 4'hF;
    W_A[84][15] = 4'hF;
    W_A[85][15] = 4'hC;
    W_A[86][15] = 4'hC;
    W_A[87][15] = 4'hC;
    W_A[88][15] = 4'hD;
    W_A[89][15] = 4'hF;
    W_A[90][15] = 4'hF;
    W_A[91][15] = 4'hD;
    W_A[92][15] = 4'hC;
    W_A[93][15] = 4'hC;
    W_A[94][15] = 4'hC;
    W_A[95][15] = 4'hF;
    W_A[96][15] = 4'hF;
    W_A[97][15] = 4'hF;
    W_A[98][15] = 4'hF;
    W_A[99][15] = 4'hF;
    W_A[100][15] = 4'hF;
    W_A[101][15] = 4'hF;
    W_A[102][15] = 4'hC;
    W_A[103][15] = 4'hC;
    W_A[104][15] = 4'hC;
    W_A[105][15] = 4'hD;
    W_A[106][15] = 4'hF;
    W_A[107][15] = 4'hF;
    W_A[0][16] = 4'hF;
    W_A[1][16] = 4'hF;
    W_A[2][16] = 4'hE;
    W_A[3][16] = 4'hD;
    W_A[4][16] = 4'hD;
    W_A[5][16] = 4'hD;
    W_A[6][16] = 4'hD;
    W_A[7][16] = 4'hD;
    W_A[8][16] = 4'hD;
    W_A[9][16] = 4'hD;
    W_A[10][16] = 4'hD;
    W_A[11][16] = 4'hD;
    W_A[12][16] = 4'hD;
    W_A[13][16] = 4'hD;
    W_A[14][16] = 4'hD;
    W_A[15][16] = 4'hD;
    W_A[16][16] = 4'hD;
    W_A[17][16] = 4'hD;
    W_A[18][16] = 4'hD;
    W_A[19][16] = 4'hD;
    W_A[20][16] = 4'hF;
    W_A[21][16] = 4'hF;
    W_A[22][16] = 4'hF;
    W_A[23][16] = 4'hD;
    W_A[24][16] = 4'hC;
    W_A[25][16] = 4'hC;
    W_A[26][16] = 4'hC;
    W_A[27][16] = 4'hC;
    W_A[28][16] = 4'hC;
    W_A[29][16] = 4'hC;
    W_A[30][16] = 4'hD;
    W_A[31][16] = 4'hF;
    W_A[32][16] = 4'hF;
    W_A[33][16] = 4'hF;
    W_A[34][16] = 4'hF;
    W_A[35][16] = 4'hF;
    W_A[36][16] = 4'hF;
    W_A[37][16] = 4'hF;
    W_A[38][16] = 4'hF;
    W_A[39][16] = 4'hF;
    W_A[40][16] = 4'hF;
    W_A[41][16] = 4'hF;
    W_A[42][16] = 4'hF;
    W_A[43][16] = 4'hF;
    W_A[44][16] = 4'hC;
    W_A[45][16] = 4'hC;
    W_A[46][16] = 4'hC;
    W_A[47][16] = 4'hC;
    W_A[48][16] = 4'hC;
    W_A[49][16] = 4'hC;
    W_A[50][16] = 4'hC;
    W_A[51][16] = 4'hC;
    W_A[52][16] = 4'hC;
    W_A[53][16] = 4'hC;
    W_A[54][16] = 4'hD;
    W_A[55][16] = 4'hF;
    W_A[56][16] = 4'hF;
    W_A[57][16] = 4'hD;
    W_A[58][16] = 4'hC;
    W_A[59][16] = 4'hC;
    W_A[60][16] = 4'hC;
    W_A[61][16] = 4'hC;
    W_A[62][16] = 4'hC;
    W_A[63][16] = 4'hC;
    W_A[64][16] = 4'hC;
    W_A[65][16] = 4'hC;
    W_A[66][16] = 4'hC;
    W_A[67][16] = 4'hC;
    W_A[68][16] = 4'hF;
    W_A[69][16] = 4'hF;
    W_A[70][16] = 4'hF;
    W_A[71][16] = 4'hF;
    W_A[72][16] = 4'hF;
    W_A[73][16] = 4'hF;
    W_A[74][16] = 4'hF;
    W_A[75][16] = 4'hF;
    W_A[76][16] = 4'hF;
    W_A[77][16] = 4'hF;
    W_A[78][16] = 4'hC;
    W_A[79][16] = 4'hC;
    W_A[80][16] = 4'hC;
    W_A[81][16] = 4'hC;
    W_A[82][16] = 4'hC;
    W_A[83][16] = 4'hC;
    W_A[84][16] = 4'hC;
    W_A[85][16] = 4'hF;
    W_A[86][16] = 4'hF;
    W_A[87][16] = 4'hF;
    W_A[88][16] = 4'hF;
    W_A[89][16] = 4'hF;
    W_A[90][16] = 4'hF;
    W_A[91][16] = 4'hD;
    W_A[92][16] = 4'hC;
    W_A[93][16] = 4'hC;
    W_A[94][16] = 4'hC;
    W_A[95][16] = 4'hF;
    W_A[96][16] = 4'hF;
    W_A[97][16] = 4'hF;
    W_A[98][16] = 4'hF;
    W_A[99][16] = 4'hF;
    W_A[100][16] = 4'hF;
    W_A[101][16] = 4'hF;
    W_A[102][16] = 4'hC;
    W_A[103][16] = 4'hC;
    W_A[104][16] = 4'hC;
    W_A[105][16] = 4'hD;
    W_A[106][16] = 4'hF;
    W_A[107][16] = 4'hF;
    W_A[0][17] = 4'hF;
    W_A[1][17] = 4'hF;
    W_A[2][17] = 4'hF;
    W_A[3][17] = 4'hF;
    W_A[4][17] = 4'hF;
    W_A[5][17] = 4'hF;
    W_A[6][17] = 4'hC;
    W_A[7][17] = 4'hC;
    W_A[8][17] = 4'hC;
    W_A[9][17] = 4'hD;
    W_A[10][17] = 4'hF;
    W_A[11][17] = 4'hF;
    W_A[12][17] = 4'hF;
    W_A[13][17] = 4'hC;
    W_A[14][17] = 4'hC;
    W_A[15][17] = 4'hC;
    W_A[16][17] = 4'hD;
    W_A[17][17] = 4'hF;
    W_A[18][17] = 4'hF;
    W_A[19][17] = 4'hF;
    W_A[20][17] = 4'hF;
    W_A[21][17] = 4'hF;
    W_A[22][17] = 4'hF;
    W_A[23][17] = 4'hF;
    W_A[24][17] = 4'hF;
    W_A[25][17] = 4'hF;
    W_A[26][17] = 4'hF;
    W_A[27][17] = 4'hC;
    W_A[28][17] = 4'hC;
    W_A[29][17] = 4'hC;
    W_A[30][17] = 4'hC;
    W_A[31][17] = 4'hC;
    W_A[32][17] = 4'hC;
    W_A[33][17] = 4'hC;
    W_A[34][17] = 4'hF;
    W_A[35][17] = 4'hF;
    W_A[36][17] = 4'hF;
    W_A[37][17] = 4'hF;
    W_A[38][17] = 4'hF;
    W_A[39][17] = 4'hF;
    W_A[40][17] = 4'hF;
    W_A[41][17] = 4'hF;
    W_A[42][17] = 4'hF;
    W_A[43][17] = 4'hF;
    W_A[44][17] = 4'hC;
    W_A[45][17] = 4'hC;
    W_A[46][17] = 4'hC;
    W_A[47][17] = 4'hC;
    W_A[48][17] = 4'hC;
    W_A[49][17] = 4'hC;
    W_A[50][17] = 4'hC;
    W_A[51][17] = 4'hC;
    W_A[52][17] = 4'hC;
    W_A[53][17] = 4'hC;
    W_A[54][17] = 4'hD;
    W_A[55][17] = 4'hF;
    W_A[56][17] = 4'hF;
    W_A[57][17] = 4'hD;
    W_A[58][17] = 4'hC;
    W_A[59][17] = 4'hC;
    W_A[60][17] = 4'hC;
    W_A[61][17] = 4'hC;
    W_A[62][17] = 4'hC;
    W_A[63][17] = 4'hC;
    W_A[64][17] = 4'hC;
    W_A[65][17] = 4'hC;
    W_A[66][17] = 4'hC;
    W_A[67][17] = 4'hC;
    W_A[68][17] = 4'hF;
    W_A[69][17] = 4'hF;
    W_A[70][17] = 4'hF;
    W_A[71][17] = 4'hF;
    W_A[72][17] = 4'hF;
    W_A[73][17] = 4'hF;
    W_A[74][17] = 4'hF;
    W_A[75][17] = 4'hF;
    W_A[76][17] = 4'hF;
    W_A[77][17] = 4'hF;
    W_A[78][17] = 4'hC;
    W_A[79][17] = 4'hC;
    W_A[80][17] = 4'hC;
    W_A[81][17] = 4'hC;
    W_A[82][17] = 4'hC;
    W_A[83][17] = 4'hC;
    W_A[84][17] = 4'hC;
    W_A[85][17] = 4'hF;
    W_A[86][17] = 4'hF;
    W_A[87][17] = 4'hF;
    W_A[88][17] = 4'hF;
    W_A[89][17] = 4'hF;
    W_A[90][17] = 4'hF;
    W_A[91][17] = 4'hD;
    W_A[92][17] = 4'hC;
    W_A[93][17] = 4'hC;
    W_A[94][17] = 4'hC;
    W_A[95][17] = 4'hF;
    W_A[96][17] = 4'hF;
    W_A[97][17] = 4'hF;
    W_A[98][17] = 4'hF;
    W_A[99][17] = 4'hF;
    W_A[100][17] = 4'hF;
    W_A[101][17] = 4'hF;
    W_A[102][17] = 4'hC;
    W_A[103][17] = 4'hC;
    W_A[104][17] = 4'hC;
    W_A[105][17] = 4'hD;
    W_A[106][17] = 4'hF;
    W_A[107][17] = 4'hF;
    W_A[0][18] = 4'hF;
    W_A[1][18] = 4'hF;
    W_A[2][18] = 4'hF;
    W_A[3][18] = 4'hF;
    W_A[4][18] = 4'hF;
    W_A[5][18] = 4'hF;
    W_A[6][18] = 4'hC;
    W_A[7][18] = 4'hC;
    W_A[8][18] = 4'hC;
    W_A[9][18] = 4'hD;
    W_A[10][18] = 4'hF;
    W_A[11][18] = 4'hF;
    W_A[12][18] = 4'hF;
    W_A[13][18] = 4'hC;
    W_A[14][18] = 4'hC;
    W_A[15][18] = 4'hC;
    W_A[16][18] = 4'hD;
    W_A[17][18] = 4'hF;
    W_A[18][18] = 4'hF;
    W_A[19][18] = 4'hF;
    W_A[20][18] = 4'hF;
    W_A[21][18] = 4'hF;
    W_A[22][18] = 4'hF;
    W_A[23][18] = 4'hF;
    W_A[24][18] = 4'hF;
    W_A[25][18] = 4'hF;
    W_A[26][18] = 4'hF;
    W_A[27][18] = 4'hC;
    W_A[28][18] = 4'hC;
    W_A[29][18] = 4'hC;
    W_A[30][18] = 4'hC;
    W_A[31][18] = 4'hC;
    W_A[32][18] = 4'hC;
    W_A[33][18] = 4'hC;
    W_A[34][18] = 4'hF;
    W_A[35][18] = 4'hF;
    W_A[36][18] = 4'hF;
    W_A[37][18] = 4'hF;
    W_A[38][18] = 4'hF;
    W_A[39][18] = 4'hF;
    W_A[40][18] = 4'hF;
    W_A[41][18] = 4'hF;
    W_A[42][18] = 4'hF;
    W_A[43][18] = 4'hF;
    W_A[44][18] = 4'hC;
    W_A[45][18] = 4'hC;
    W_A[46][18] = 4'hC;
    W_A[47][18] = 4'hC;
    W_A[48][18] = 4'hC;
    W_A[49][18] = 4'hC;
    W_A[50][18] = 4'hC;
    W_A[51][18] = 4'hC;
    W_A[52][18] = 4'hC;
    W_A[53][18] = 4'hC;
    W_A[54][18] = 4'hD;
    W_A[55][18] = 4'hF;
    W_A[56][18] = 4'hF;
    W_A[57][18] = 4'hD;
    W_A[58][18] = 4'hC;
    W_A[59][18] = 4'hC;
    W_A[60][18] = 4'hC;
    W_A[61][18] = 4'hC;
    W_A[62][18] = 4'hC;
    W_A[63][18] = 4'hC;
    W_A[64][18] = 4'hC;
    W_A[65][18] = 4'hC;
    W_A[66][18] = 4'hC;
    W_A[67][18] = 4'hC;
    W_A[68][18] = 4'hF;
    W_A[69][18] = 4'hF;
    W_A[70][18] = 4'hF;
    W_A[71][18] = 4'hF;
    W_A[72][18] = 4'hF;
    W_A[73][18] = 4'hF;
    W_A[74][18] = 4'hF;
    W_A[75][18] = 4'hF;
    W_A[76][18] = 4'hF;
    W_A[77][18] = 4'hF;
    W_A[78][18] = 4'hC;
    W_A[79][18] = 4'hC;
    W_A[80][18] = 4'hC;
    W_A[81][18] = 4'hC;
    W_A[82][18] = 4'hC;
    W_A[83][18] = 4'hC;
    W_A[84][18] = 4'hC;
    W_A[85][18] = 4'hF;
    W_A[86][18] = 4'hF;
    W_A[87][18] = 4'hF;
    W_A[88][18] = 4'hF;
    W_A[89][18] = 4'hF;
    W_A[90][18] = 4'hF;
    W_A[91][18] = 4'hD;
    W_A[92][18] = 4'hC;
    W_A[93][18] = 4'hC;
    W_A[94][18] = 4'hC;
    W_A[95][18] = 4'hF;
    W_A[96][18] = 4'hF;
    W_A[97][18] = 4'hF;
    W_A[98][18] = 4'hF;
    W_A[99][18] = 4'hF;
    W_A[100][18] = 4'hF;
    W_A[101][18] = 4'hF;
    W_A[102][18] = 4'hC;
    W_A[103][18] = 4'hC;
    W_A[104][18] = 4'hC;
    W_A[105][18] = 4'hD;
    W_A[106][18] = 4'hF;
    W_A[107][18] = 4'hF;
    W_A[0][19] = 4'hF;
    W_A[1][19] = 4'hF;
    W_A[2][19] = 4'hF;
    W_A[3][19] = 4'hF;
    W_A[4][19] = 4'hF;
    W_A[5][19] = 4'hF;
    W_A[6][19] = 4'hC;
    W_A[7][19] = 4'hC;
    W_A[8][19] = 4'hC;
    W_A[9][19] = 4'hD;
    W_A[10][19] = 4'hF;
    W_A[11][19] = 4'hF;
    W_A[12][19] = 4'hF;
    W_A[13][19] = 4'hC;
    W_A[14][19] = 4'hC;
    W_A[15][19] = 4'hC;
    W_A[16][19] = 4'hD;
    W_A[17][19] = 4'hF;
    W_A[18][19] = 4'hF;
    W_A[19][19] = 4'hF;
    W_A[20][19] = 4'hF;
    W_A[21][19] = 4'hF;
    W_A[22][19] = 4'hF;
    W_A[23][19] = 4'hF;
    W_A[24][19] = 4'hF;
    W_A[25][19] = 4'hF;
    W_A[26][19] = 4'hF;
    W_A[27][19] = 4'hC;
    W_A[28][19] = 4'hC;
    W_A[29][19] = 4'hC;
    W_A[30][19] = 4'hC;
    W_A[31][19] = 4'hC;
    W_A[32][19] = 4'hC;
    W_A[33][19] = 4'hC;
    W_A[34][19] = 4'hF;
    W_A[35][19] = 4'hF;
    W_A[36][19] = 4'hF;
    W_A[37][19] = 4'hF;
    W_A[38][19] = 4'hF;
    W_A[39][19] = 4'hF;
    W_A[40][19] = 4'hF;
    W_A[41][19] = 4'hF;
    W_A[42][19] = 4'hF;
    W_A[43][19] = 4'hF;
    W_A[44][19] = 4'hC;
    W_A[45][19] = 4'hC;
    W_A[46][19] = 4'hC;
    W_A[47][19] = 4'hC;
    W_A[48][19] = 4'hC;
    W_A[49][19] = 4'hC;
    W_A[50][19] = 4'hC;
    W_A[51][19] = 4'hC;
    W_A[52][19] = 4'hC;
    W_A[53][19] = 4'hC;
    W_A[54][19] = 4'hD;
    W_A[55][19] = 4'hF;
    W_A[56][19] = 4'hF;
    W_A[57][19] = 4'hD;
    W_A[58][19] = 4'hC;
    W_A[59][19] = 4'hC;
    W_A[60][19] = 4'hC;
    W_A[61][19] = 4'hC;
    W_A[62][19] = 4'hC;
    W_A[63][19] = 4'hC;
    W_A[64][19] = 4'hC;
    W_A[65][19] = 4'hC;
    W_A[66][19] = 4'hC;
    W_A[67][19] = 4'hC;
    W_A[68][19] = 4'hF;
    W_A[69][19] = 4'hF;
    W_A[70][19] = 4'hF;
    W_A[71][19] = 4'hF;
    W_A[72][19] = 4'hF;
    W_A[73][19] = 4'hF;
    W_A[74][19] = 4'hF;
    W_A[75][19] = 4'hF;
    W_A[76][19] = 4'hF;
    W_A[77][19] = 4'hF;
    W_A[78][19] = 4'hC;
    W_A[79][19] = 4'hC;
    W_A[80][19] = 4'hC;
    W_A[81][19] = 4'hC;
    W_A[82][19] = 4'hC;
    W_A[83][19] = 4'hC;
    W_A[84][19] = 4'hC;
    W_A[85][19] = 4'hF;
    W_A[86][19] = 4'hF;
    W_A[87][19] = 4'hF;
    W_A[88][19] = 4'hF;
    W_A[89][19] = 4'hF;
    W_A[90][19] = 4'hF;
    W_A[91][19] = 4'hD;
    W_A[92][19] = 4'hC;
    W_A[93][19] = 4'hC;
    W_A[94][19] = 4'hC;
    W_A[95][19] = 4'hF;
    W_A[96][19] = 4'hF;
    W_A[97][19] = 4'hF;
    W_A[98][19] = 4'hF;
    W_A[99][19] = 4'hF;
    W_A[100][19] = 4'hF;
    W_A[101][19] = 4'hF;
    W_A[102][19] = 4'hC;
    W_A[103][19] = 4'hC;
    W_A[104][19] = 4'hC;
    W_A[105][19] = 4'hD;
    W_A[106][19] = 4'hF;
    W_A[107][19] = 4'hF;
    W_A[0][20] = 4'hF;
    W_A[1][20] = 4'hF;
    W_A[2][20] = 4'hF;
    W_A[3][20] = 4'hF;
    W_A[4][20] = 4'hF;
    W_A[5][20] = 4'hF;
    W_A[6][20] = 4'hF;
    W_A[7][20] = 4'hF;
    W_A[8][20] = 4'hF;
    W_A[9][20] = 4'hF;
    W_A[10][20] = 4'hF;
    W_A[11][20] = 4'hF;
    W_A[12][20] = 4'hF;
    W_A[13][20] = 4'hF;
    W_A[14][20] = 4'hF;
    W_A[15][20] = 4'hF;
    W_A[16][20] = 4'hF;
    W_A[17][20] = 4'hF;
    W_A[18][20] = 4'hF;
    W_A[19][20] = 4'hF;
    W_A[20][20] = 4'hF;
    W_A[21][20] = 4'hF;
    W_A[22][20] = 4'hF;
    W_A[23][20] = 4'hF;
    W_A[24][20] = 4'hF;
    W_A[25][20] = 4'hF;
    W_A[26][20] = 4'hF;
    W_A[27][20] = 4'hF;
    W_A[28][20] = 4'hF;
    W_A[29][20] = 4'hF;
    W_A[30][20] = 4'hF;
    W_A[31][20] = 4'hF;
    W_A[32][20] = 4'hF;
    W_A[33][20] = 4'hF;
    W_A[34][20] = 4'hF;
    W_A[35][20] = 4'hF;
    W_A[36][20] = 4'hF;
    W_A[37][20] = 4'hF;
    W_A[38][20] = 4'hF;
    W_A[39][20] = 4'hF;
    W_A[40][20] = 4'hF;
    W_A[41][20] = 4'hF;
    W_A[42][20] = 4'hF;
    W_A[43][20] = 4'hF;
    W_A[44][20] = 4'hF;
    W_A[45][20] = 4'hF;
    W_A[46][20] = 4'hF;
    W_A[47][20] = 4'hF;
    W_A[48][20] = 4'hF;
    W_A[49][20] = 4'hF;
    W_A[50][20] = 4'hF;
    W_A[51][20] = 4'hF;
    W_A[52][20] = 4'hF;
    W_A[53][20] = 4'hF;
    W_A[54][20] = 4'hF;
    W_A[55][20] = 4'hF;
    W_A[56][20] = 4'hF;
    W_A[57][20] = 4'hD;
    W_A[58][20] = 4'hC;
    W_A[59][20] = 4'hC;
    W_A[60][20] = 4'hC;
    W_A[61][20] = 4'hF;
    W_A[62][20] = 4'hF;
    W_A[63][20] = 4'hF;
    W_A[64][20] = 4'hF;
    W_A[65][20] = 4'hF;
    W_A[66][20] = 4'hF;
    W_A[67][20] = 4'hF;
    W_A[68][20] = 4'hF;
    W_A[69][20] = 4'hF;
    W_A[70][20] = 4'hF;
    W_A[71][20] = 4'hF;
    W_A[72][20] = 4'hF;
    W_A[73][20] = 4'hF;
    W_A[74][20] = 4'hF;
    W_A[75][20] = 4'hF;
    W_A[76][20] = 4'hF;
    W_A[77][20] = 4'hF;
    W_A[78][20] = 4'hF;
    W_A[79][20] = 4'hF;
    W_A[80][20] = 4'hF;
    W_A[81][20] = 4'hF;
    W_A[82][20] = 4'hF;
    W_A[83][20] = 4'hF;
    W_A[84][20] = 4'hF;
    W_A[85][20] = 4'hF;
    W_A[86][20] = 4'hF;
    W_A[87][20] = 4'hF;
    W_A[88][20] = 4'hF;
    W_A[89][20] = 4'hF;
    W_A[90][20] = 4'hF;
    W_A[91][20] = 4'hF;
    W_A[92][20] = 4'hF;
    W_A[93][20] = 4'hF;
    W_A[94][20] = 4'hF;
    W_A[95][20] = 4'hF;
    W_A[96][20] = 4'hF;
    W_A[97][20] = 4'hF;
    W_A[98][20] = 4'hF;
    W_A[99][20] = 4'hF;
    W_A[100][20] = 4'hF;
    W_A[101][20] = 4'hF;
    W_A[102][20] = 4'hF;
    W_A[103][20] = 4'hF;
    W_A[104][20] = 4'hF;
    W_A[105][20] = 4'hF;
    W_A[106][20] = 4'hF;
    W_A[107][20] = 4'hF;
    W_A[0][21] = 4'hF;
    W_A[1][21] = 4'hF;
    W_A[2][21] = 4'hF;
    W_A[3][21] = 4'hF;
    W_A[4][21] = 4'hF;
    W_A[5][21] = 4'hF;
    W_A[6][21] = 4'hF;
    W_A[7][21] = 4'hF;
    W_A[8][21] = 4'hF;
    W_A[9][21] = 4'hF;
    W_A[10][21] = 4'hF;
    W_A[11][21] = 4'hF;
    W_A[12][21] = 4'hF;
    W_A[13][21] = 4'hF;
    W_A[14][21] = 4'hF;
    W_A[15][21] = 4'hF;
    W_A[16][21] = 4'hF;
    W_A[17][21] = 4'hF;
    W_A[18][21] = 4'hF;
    W_A[19][21] = 4'hF;
    W_A[20][21] = 4'hF;
    W_A[21][21] = 4'hF;
    W_A[22][21] = 4'hF;
    W_A[23][21] = 4'hF;
    W_A[24][21] = 4'hF;
    W_A[25][21] = 4'hF;
    W_A[26][21] = 4'hF;
    W_A[27][21] = 4'hF;
    W_A[28][21] = 4'hF;
    W_A[29][21] = 4'hF;
    W_A[30][21] = 4'hF;
    W_A[31][21] = 4'hF;
    W_A[32][21] = 4'hF;
    W_A[33][21] = 4'hF;
    W_A[34][21] = 4'hF;
    W_A[35][21] = 4'hF;
    W_A[36][21] = 4'hF;
    W_A[37][21] = 4'hF;
    W_A[38][21] = 4'hF;
    W_A[39][21] = 4'hF;
    W_A[40][21] = 4'hF;
    W_A[41][21] = 4'hF;
    W_A[42][21] = 4'hF;
    W_A[43][21] = 4'hF;
    W_A[44][21] = 4'hF;
    W_A[45][21] = 4'hF;
    W_A[46][21] = 4'hF;
    W_A[47][21] = 4'hF;
    W_A[48][21] = 4'hF;
    W_A[49][21] = 4'hF;
    W_A[50][21] = 4'hF;
    W_A[51][21] = 4'hF;
    W_A[52][21] = 4'hF;
    W_A[53][21] = 4'hF;
    W_A[54][21] = 4'hF;
    W_A[55][21] = 4'hF;
    W_A[56][21] = 4'hF;
    W_A[57][21] = 4'hD;
    W_A[58][21] = 4'hC;
    W_A[59][21] = 4'hC;
    W_A[60][21] = 4'hC;
    W_A[61][21] = 4'hF;
    W_A[62][21] = 4'hF;
    W_A[63][21] = 4'hF;
    W_A[64][21] = 4'hF;
    W_A[65][21] = 4'hF;
    W_A[66][21] = 4'hF;
    W_A[67][21] = 4'hF;
    W_A[68][21] = 4'hF;
    W_A[69][21] = 4'hF;
    W_A[70][21] = 4'hF;
    W_A[71][21] = 4'hF;
    W_A[72][21] = 4'hF;
    W_A[73][21] = 4'hF;
    W_A[74][21] = 4'hF;
    W_A[75][21] = 4'hF;
    W_A[76][21] = 4'hF;
    W_A[77][21] = 4'hF;
    W_A[78][21] = 4'hF;
    W_A[79][21] = 4'hF;
    W_A[80][21] = 4'hF;
    W_A[81][21] = 4'hF;
    W_A[82][21] = 4'hF;
    W_A[83][21] = 4'hF;
    W_A[84][21] = 4'hF;
    W_A[85][21] = 4'hF;
    W_A[86][21] = 4'hF;
    W_A[87][21] = 4'hF;
    W_A[88][21] = 4'hF;
    W_A[89][21] = 4'hF;
    W_A[90][21] = 4'hF;
    W_A[91][21] = 4'hF;
    W_A[92][21] = 4'hF;
    W_A[93][21] = 4'hF;
    W_A[94][21] = 4'hF;
    W_A[95][21] = 4'hF;
    W_A[96][21] = 4'hF;
    W_A[97][21] = 4'hF;
    W_A[98][21] = 4'hF;
    W_A[99][21] = 4'hF;
    W_A[100][21] = 4'hF;
    W_A[101][21] = 4'hF;
    W_A[102][21] = 4'hF;
    W_A[103][21] = 4'hF;
    W_A[104][21] = 4'hF;
    W_A[105][21] = 4'hF;
    W_A[106][21] = 4'hF;
    W_A[107][21] = 4'hF;
    W_A[0][22] = 4'hF;
    W_A[1][22] = 4'hF;
    W_A[2][22] = 4'hF;
    W_A[3][22] = 4'hF;
    W_A[4][22] = 4'hF;
    W_A[5][22] = 4'hF;
    W_A[6][22] = 4'hF;
    W_A[7][22] = 4'hF;
    W_A[8][22] = 4'hF;
    W_A[9][22] = 4'hF;
    W_A[10][22] = 4'hF;
    W_A[11][22] = 4'hF;
    W_A[12][22] = 4'hF;
    W_A[13][22] = 4'hF;
    W_A[14][22] = 4'hF;
    W_A[15][22] = 4'hF;
    W_A[16][22] = 4'hF;
    W_A[17][22] = 4'hF;
    W_A[18][22] = 4'hF;
    W_A[19][22] = 4'hF;
    W_A[20][22] = 4'hF;
    W_A[21][22] = 4'hF;
    W_A[22][22] = 4'hF;
    W_A[23][22] = 4'hF;
    W_A[24][22] = 4'hF;
    W_A[25][22] = 4'hF;
    W_A[26][22] = 4'hF;
    W_A[27][22] = 4'hF;
    W_A[28][22] = 4'hF;
    W_A[29][22] = 4'hF;
    W_A[30][22] = 4'hF;
    W_A[31][22] = 4'hF;
    W_A[32][22] = 4'hF;
    W_A[33][22] = 4'hF;
    W_A[34][22] = 4'hF;
    W_A[35][22] = 4'hF;
    W_A[36][22] = 4'hF;
    W_A[37][22] = 4'hF;
    W_A[38][22] = 4'hF;
    W_A[39][22] = 4'hF;
    W_A[40][22] = 4'hF;
    W_A[41][22] = 4'hF;
    W_A[42][22] = 4'hF;
    W_A[43][22] = 4'hF;
    W_A[44][22] = 4'hF;
    W_A[45][22] = 4'hF;
    W_A[46][22] = 4'hF;
    W_A[47][22] = 4'hF;
    W_A[48][22] = 4'hF;
    W_A[49][22] = 4'hF;
    W_A[50][22] = 4'hF;
    W_A[51][22] = 4'hF;
    W_A[52][22] = 4'hF;
    W_A[53][22] = 4'hF;
    W_A[54][22] = 4'hF;
    W_A[55][22] = 4'hF;
    W_A[56][22] = 4'hF;
    W_A[57][22] = 4'hD;
    W_A[58][22] = 4'hC;
    W_A[59][22] = 4'hC;
    W_A[60][22] = 4'hC;
    W_A[61][22] = 4'hF;
    W_A[62][22] = 4'hF;
    W_A[63][22] = 4'hF;
    W_A[64][22] = 4'hF;
    W_A[65][22] = 4'hF;
    W_A[66][22] = 4'hF;
    W_A[67][22] = 4'hF;
    W_A[68][22] = 4'hF;
    W_A[69][22] = 4'hF;
    W_A[70][22] = 4'hF;
    W_A[71][22] = 4'hF;
    W_A[72][22] = 4'hF;
    W_A[73][22] = 4'hF;
    W_A[74][22] = 4'hF;
    W_A[75][22] = 4'hF;
    W_A[76][22] = 4'hF;
    W_A[77][22] = 4'hF;
    W_A[78][22] = 4'hF;
    W_A[79][22] = 4'hF;
    W_A[80][22] = 4'hF;
    W_A[81][22] = 4'hF;
    W_A[82][22] = 4'hF;
    W_A[83][22] = 4'hF;
    W_A[84][22] = 4'hF;
    W_A[85][22] = 4'hF;
    W_A[86][22] = 4'hF;
    W_A[87][22] = 4'hF;
    W_A[88][22] = 4'hF;
    W_A[89][22] = 4'hF;
    W_A[90][22] = 4'hF;
    W_A[91][22] = 4'hF;
    W_A[92][22] = 4'hF;
    W_A[93][22] = 4'hF;
    W_A[94][22] = 4'hF;
    W_A[95][22] = 4'hF;
    W_A[96][22] = 4'hF;
    W_A[97][22] = 4'hF;
    W_A[98][22] = 4'hF;
    W_A[99][22] = 4'hF;
    W_A[100][22] = 4'hF;
    W_A[101][22] = 4'hF;
    W_A[102][22] = 4'hF;
    W_A[103][22] = 4'hF;
    W_A[104][22] = 4'hF;
    W_A[105][22] = 4'hF;
    W_A[106][22] = 4'hF;
    W_A[107][22] = 4'hF;
    W_A[0][23] = 4'hF;
    W_A[1][23] = 4'hF;
    W_A[2][23] = 4'hF;
    W_A[3][23] = 4'hF;
    W_A[4][23] = 4'hF;
    W_A[5][23] = 4'hF;
    W_A[6][23] = 4'hF;
    W_A[7][23] = 4'hF;
    W_A[8][23] = 4'hF;
    W_A[9][23] = 4'hF;
    W_A[10][23] = 4'hF;
    W_A[11][23] = 4'hF;
    W_A[12][23] = 4'hF;
    W_A[13][23] = 4'hF;
    W_A[14][23] = 4'hF;
    W_A[15][23] = 4'hF;
    W_A[16][23] = 4'hF;
    W_A[17][23] = 4'hF;
    W_A[18][23] = 4'hF;
    W_A[19][23] = 4'hF;
    W_A[20][23] = 4'hF;
    W_A[21][23] = 4'hF;
    W_A[22][23] = 4'hF;
    W_A[23][23] = 4'hF;
    W_A[24][23] = 4'hF;
    W_A[25][23] = 4'hF;
    W_A[26][23] = 4'hF;
    W_A[27][23] = 4'hF;
    W_A[28][23] = 4'hF;
    W_A[29][23] = 4'hF;
    W_A[30][23] = 4'hF;
    W_A[31][23] = 4'hF;
    W_A[32][23] = 4'hF;
    W_A[33][23] = 4'hF;
    W_A[34][23] = 4'hF;
    W_A[35][23] = 4'hF;
    W_A[36][23] = 4'hF;
    W_A[37][23] = 4'hF;
    W_A[38][23] = 4'hF;
    W_A[39][23] = 4'hF;
    W_A[40][23] = 4'hF;
    W_A[41][23] = 4'hF;
    W_A[42][23] = 4'hF;
    W_A[43][23] = 4'hF;
    W_A[44][23] = 4'hF;
    W_A[45][23] = 4'hF;
    W_A[46][23] = 4'hF;
    W_A[47][23] = 4'hF;
    W_A[48][23] = 4'hF;
    W_A[49][23] = 4'hF;
    W_A[50][23] = 4'hF;
    W_A[51][23] = 4'hF;
    W_A[52][23] = 4'hF;
    W_A[53][23] = 4'hF;
    W_A[54][23] = 4'hF;
    W_A[55][23] = 4'hF;
    W_A[56][23] = 4'hF;
    W_A[57][23] = 4'hD;
    W_A[58][23] = 4'hC;
    W_A[59][23] = 4'hC;
    W_A[60][23] = 4'hC;
    W_A[61][23] = 4'hF;
    W_A[62][23] = 4'hF;
    W_A[63][23] = 4'hF;
    W_A[64][23] = 4'hF;
    W_A[65][23] = 4'hF;
    W_A[66][23] = 4'hF;
    W_A[67][23] = 4'hF;
    W_A[68][23] = 4'hF;
    W_A[69][23] = 4'hF;
    W_A[70][23] = 4'hF;
    W_A[71][23] = 4'hF;
    W_A[72][23] = 4'hF;
    W_A[73][23] = 4'hF;
    W_A[74][23] = 4'hF;
    W_A[75][23] = 4'hF;
    W_A[76][23] = 4'hF;
    W_A[77][23] = 4'hF;
    W_A[78][23] = 4'hF;
    W_A[79][23] = 4'hF;
    W_A[80][23] = 4'hF;
    W_A[81][23] = 4'hF;
    W_A[82][23] = 4'hF;
    W_A[83][23] = 4'hF;
    W_A[84][23] = 4'hF;
    W_A[85][23] = 4'hF;
    W_A[86][23] = 4'hF;
    W_A[87][23] = 4'hF;
    W_A[88][23] = 4'hF;
    W_A[89][23] = 4'hF;
    W_A[90][23] = 4'hF;
    W_A[91][23] = 4'hF;
    W_A[92][23] = 4'hF;
    W_A[93][23] = 4'hF;
    W_A[94][23] = 4'hF;
    W_A[95][23] = 4'hF;
    W_A[96][23] = 4'hF;
    W_A[97][23] = 4'hF;
    W_A[98][23] = 4'hF;
    W_A[99][23] = 4'hF;
    W_A[100][23] = 4'hF;
    W_A[101][23] = 4'hF;
    W_A[102][23] = 4'hF;
    W_A[103][23] = 4'hF;
    W_A[104][23] = 4'hF;
    W_A[105][23] = 4'hF;
    W_A[106][23] = 4'hF;
    W_A[107][23] = 4'hF;
    W_A[0][24] = 4'hF;
    W_A[1][24] = 4'hF;
    W_A[2][24] = 4'hF;
    W_A[3][24] = 4'hF;
    W_A[4][24] = 4'hF;
    W_A[5][24] = 4'hF;
    W_A[6][24] = 4'hF;
    W_A[7][24] = 4'hF;
    W_A[8][24] = 4'hF;
    W_A[9][24] = 4'hF;
    W_A[10][24] = 4'hF;
    W_A[11][24] = 4'hF;
    W_A[12][24] = 4'hF;
    W_A[13][24] = 4'hF;
    W_A[14][24] = 4'hF;
    W_A[15][24] = 4'hF;
    W_A[16][24] = 4'hF;
    W_A[17][24] = 4'hF;
    W_A[18][24] = 4'hF;
    W_A[19][24] = 4'hF;
    W_A[20][24] = 4'hF;
    W_A[21][24] = 4'hF;
    W_A[22][24] = 4'hF;
    W_A[23][24] = 4'hF;
    W_A[24][24] = 4'hF;
    W_A[25][24] = 4'hF;
    W_A[26][24] = 4'hF;
    W_A[27][24] = 4'hF;
    W_A[28][24] = 4'hF;
    W_A[29][24] = 4'hF;
    W_A[30][24] = 4'hF;
    W_A[31][24] = 4'hF;
    W_A[32][24] = 4'hF;
    W_A[33][24] = 4'hF;
    W_A[34][24] = 4'hF;
    W_A[35][24] = 4'hF;
    W_A[36][24] = 4'hF;
    W_A[37][24] = 4'hF;
    W_A[38][24] = 4'hF;
    W_A[39][24] = 4'hF;
    W_A[40][24] = 4'hF;
    W_A[41][24] = 4'hF;
    W_A[42][24] = 4'hF;
    W_A[43][24] = 4'hF;
    W_A[44][24] = 4'hF;
    W_A[45][24] = 4'hF;
    W_A[46][24] = 4'hF;
    W_A[47][24] = 4'hF;
    W_A[48][24] = 4'hF;
    W_A[49][24] = 4'hF;
    W_A[50][24] = 4'hF;
    W_A[51][24] = 4'hF;
    W_A[52][24] = 4'hF;
    W_A[53][24] = 4'hF;
    W_A[54][24] = 4'hF;
    W_A[55][24] = 4'hF;
    W_A[56][24] = 4'hF;
    W_A[57][24] = 4'hD;
    W_A[58][24] = 4'hC;
    W_A[59][24] = 4'hC;
    W_A[60][24] = 4'hC;
    W_A[61][24] = 4'hF;
    W_A[62][24] = 4'hF;
    W_A[63][24] = 4'hF;
    W_A[64][24] = 4'hF;
    W_A[65][24] = 4'hF;
    W_A[66][24] = 4'hF;
    W_A[67][24] = 4'hF;
    W_A[68][24] = 4'hF;
    W_A[69][24] = 4'hF;
    W_A[70][24] = 4'hF;
    W_A[71][24] = 4'hF;
    W_A[72][24] = 4'hF;
    W_A[73][24] = 4'hF;
    W_A[74][24] = 4'hF;
    W_A[75][24] = 4'hF;
    W_A[76][24] = 4'hF;
    W_A[77][24] = 4'hF;
    W_A[78][24] = 4'hF;
    W_A[79][24] = 4'hF;
    W_A[80][24] = 4'hF;
    W_A[81][24] = 4'hF;
    W_A[82][24] = 4'hF;
    W_A[83][24] = 4'hF;
    W_A[84][24] = 4'hF;
    W_A[85][24] = 4'hF;
    W_A[86][24] = 4'hF;
    W_A[87][24] = 4'hF;
    W_A[88][24] = 4'hF;
    W_A[89][24] = 4'hF;
    W_A[90][24] = 4'hF;
    W_A[91][24] = 4'hF;
    W_A[92][24] = 4'hF;
    W_A[93][24] = 4'hF;
    W_A[94][24] = 4'hF;
    W_A[95][24] = 4'hF;
    W_A[96][24] = 4'hF;
    W_A[97][24] = 4'hF;
    W_A[98][24] = 4'hF;
    W_A[99][24] = 4'hF;
    W_A[100][24] = 4'hF;
    W_A[101][24] = 4'hF;
    W_A[102][24] = 4'hF;
    W_A[103][24] = 4'hF;
    W_A[104][24] = 4'hF;
    W_A[105][24] = 4'hF;
    W_A[106][24] = 4'hF;
    W_A[107][24] = 4'hF;
    W_A[0][25] = 4'hF;
    W_A[1][25] = 4'hF;
    W_A[2][25] = 4'hF;
    W_A[3][25] = 4'hF;
    W_A[4][25] = 4'hF;
    W_A[5][25] = 4'hF;
    W_A[6][25] = 4'hF;
    W_A[7][25] = 4'hF;
    W_A[8][25] = 4'hF;
    W_A[9][25] = 4'hF;
    W_A[10][25] = 4'hF;
    W_A[11][25] = 4'hF;
    W_A[12][25] = 4'hF;
    W_A[13][25] = 4'hF;
    W_A[14][25] = 4'hF;
    W_A[15][25] = 4'hF;
    W_A[16][25] = 4'hF;
    W_A[17][25] = 4'hF;
    W_A[18][25] = 4'hF;
    W_A[19][25] = 4'hF;
    W_A[20][25] = 4'hF;
    W_A[21][25] = 4'hF;
    W_A[22][25] = 4'hF;
    W_A[23][25] = 4'hF;
    W_A[24][25] = 4'hF;
    W_A[25][25] = 4'hF;
    W_A[26][25] = 4'hF;
    W_A[27][25] = 4'hF;
    W_A[28][25] = 4'hF;
    W_A[29][25] = 4'hF;
    W_A[30][25] = 4'hF;
    W_A[31][25] = 4'hF;
    W_A[32][25] = 4'hF;
    W_A[33][25] = 4'hF;
    W_A[34][25] = 4'hF;
    W_A[35][25] = 4'hF;
    W_A[36][25] = 4'hF;
    W_A[37][25] = 4'hF;
    W_A[38][25] = 4'hF;
    W_A[39][25] = 4'hF;
    W_A[40][25] = 4'hF;
    W_A[41][25] = 4'hF;
    W_A[42][25] = 4'hF;
    W_A[43][25] = 4'hF;
    W_A[44][25] = 4'hF;
    W_A[45][25] = 4'hF;
    W_A[46][25] = 4'hF;
    W_A[47][25] = 4'hF;
    W_A[48][25] = 4'hF;
    W_A[49][25] = 4'hF;
    W_A[50][25] = 4'hF;
    W_A[51][25] = 4'hF;
    W_A[52][25] = 4'hF;
    W_A[53][25] = 4'hF;
    W_A[54][25] = 4'hF;
    W_A[55][25] = 4'hF;
    W_A[56][25] = 4'hF;
    W_A[57][25] = 4'hD;
    W_A[58][25] = 4'hC;
    W_A[59][25] = 4'hC;
    W_A[60][25] = 4'hC;
    W_A[61][25] = 4'hF;
    W_A[62][25] = 4'hF;
    W_A[63][25] = 4'hF;
    W_A[64][25] = 4'hF;
    W_A[65][25] = 4'hF;
    W_A[66][25] = 4'hF;
    W_A[67][25] = 4'hF;
    W_A[68][25] = 4'hF;
    W_A[69][25] = 4'hF;
    W_A[70][25] = 4'hF;
    W_A[71][25] = 4'hF;
    W_A[72][25] = 4'hF;
    W_A[73][25] = 4'hF;
    W_A[74][25] = 4'hF;
    W_A[75][25] = 4'hF;
    W_A[76][25] = 4'hF;
    W_A[77][25] = 4'hF;
    W_A[78][25] = 4'hF;
    W_A[79][25] = 4'hF;
    W_A[80][25] = 4'hF;
    W_A[81][25] = 4'hF;
    W_A[82][25] = 4'hF;
    W_A[83][25] = 4'hF;
    W_A[84][25] = 4'hF;
    W_A[85][25] = 4'hF;
    W_A[86][25] = 4'hF;
    W_A[87][25] = 4'hF;
    W_A[88][25] = 4'hF;
    W_A[89][25] = 4'hF;
    W_A[90][25] = 4'hF;
    W_A[91][25] = 4'hF;
    W_A[92][25] = 4'hF;
    W_A[93][25] = 4'hF;
    W_A[94][25] = 4'hF;
    W_A[95][25] = 4'hF;
    W_A[96][25] = 4'hF;
    W_A[97][25] = 4'hF;
    W_A[98][25] = 4'hF;
    W_A[99][25] = 4'hF;
    W_A[100][25] = 4'hF;
    W_A[101][25] = 4'hF;
    W_A[102][25] = 4'hF;
    W_A[103][25] = 4'hF;
    W_A[104][25] = 4'hF;
    W_A[105][25] = 4'hF;
    W_A[106][25] = 4'hF;
    W_A[107][25] = 4'hF;
    W_A[0][26] = 4'hF;
    W_A[1][26] = 4'hF;
    W_A[2][26] = 4'hF;
    W_A[3][26] = 4'hF;
    W_A[4][26] = 4'hF;
    W_A[5][26] = 4'hF;
    W_A[6][26] = 4'hF;
    W_A[7][26] = 4'hF;
    W_A[8][26] = 4'hF;
    W_A[9][26] = 4'hF;
    W_A[10][26] = 4'hF;
    W_A[11][26] = 4'hF;
    W_A[12][26] = 4'hF;
    W_A[13][26] = 4'hF;
    W_A[14][26] = 4'hF;
    W_A[15][26] = 4'hF;
    W_A[16][26] = 4'hF;
    W_A[17][26] = 4'hF;
    W_A[18][26] = 4'hF;
    W_A[19][26] = 4'hF;
    W_A[20][26] = 4'hF;
    W_A[21][26] = 4'hF;
    W_A[22][26] = 4'hF;
    W_A[23][26] = 4'hF;
    W_A[24][26] = 4'hF;
    W_A[25][26] = 4'hF;
    W_A[26][26] = 4'hF;
    W_A[27][26] = 4'hF;
    W_A[28][26] = 4'hF;
    W_A[29][26] = 4'hF;
    W_A[30][26] = 4'hF;
    W_A[31][26] = 4'hF;
    W_A[32][26] = 4'hF;
    W_A[33][26] = 4'hF;
    W_A[34][26] = 4'hF;
    W_A[35][26] = 4'hF;
    W_A[36][26] = 4'hF;
    W_A[37][26] = 4'hF;
    W_A[38][26] = 4'hF;
    W_A[39][26] = 4'hF;
    W_A[40][26] = 4'hF;
    W_A[41][26] = 4'hF;
    W_A[42][26] = 4'hF;
    W_A[43][26] = 4'hF;
    W_A[44][26] = 4'hF;
    W_A[45][26] = 4'hF;
    W_A[46][26] = 4'hF;
    W_A[47][26] = 4'hF;
    W_A[48][26] = 4'hF;
    W_A[49][26] = 4'hF;
    W_A[50][26] = 4'hF;
    W_A[51][26] = 4'hF;
    W_A[52][26] = 4'hF;
    W_A[53][26] = 4'hF;
    W_A[54][26] = 4'hF;
    W_A[55][26] = 4'hF;
    W_A[56][26] = 4'hF;
    W_A[57][26] = 4'hD;
    W_A[58][26] = 4'hC;
    W_A[59][26] = 4'hC;
    W_A[60][26] = 4'hC;
    W_A[61][26] = 4'hF;
    W_A[62][26] = 4'hF;
    W_A[63][26] = 4'hF;
    W_A[64][26] = 4'hF;
    W_A[65][26] = 4'hF;
    W_A[66][26] = 4'hF;
    W_A[67][26] = 4'hF;
    W_A[68][26] = 4'hF;
    W_A[69][26] = 4'hF;
    W_A[70][26] = 4'hF;
    W_A[71][26] = 4'hF;
    W_A[72][26] = 4'hF;
    W_A[73][26] = 4'hF;
    W_A[74][26] = 4'hF;
    W_A[75][26] = 4'hF;
    W_A[76][26] = 4'hF;
    W_A[77][26] = 4'hF;
    W_A[78][26] = 4'hF;
    W_A[79][26] = 4'hF;
    W_A[80][26] = 4'hF;
    W_A[81][26] = 4'hF;
    W_A[82][26] = 4'hF;
    W_A[83][26] = 4'hF;
    W_A[84][26] = 4'hF;
    W_A[85][26] = 4'hF;
    W_A[86][26] = 4'hF;
    W_A[87][26] = 4'hF;
    W_A[88][26] = 4'hF;
    W_A[89][26] = 4'hF;
    W_A[90][26] = 4'hF;
    W_A[91][26] = 4'hF;
    W_A[92][26] = 4'hF;
    W_A[93][26] = 4'hF;
    W_A[94][26] = 4'hF;
    W_A[95][26] = 4'hF;
    W_A[96][26] = 4'hF;
    W_A[97][26] = 4'hF;
    W_A[98][26] = 4'hF;
    W_A[99][26] = 4'hF;
    W_A[100][26] = 4'hF;
    W_A[101][26] = 4'hF;
    W_A[102][26] = 4'hF;
    W_A[103][26] = 4'hF;
    W_A[104][26] = 4'hF;
    W_A[105][26] = 4'hF;
    W_A[106][26] = 4'hF;
    W_A[107][26] = 4'hF;
    W_A[0][27] = 4'hF;
    W_A[1][27] = 4'hF;
    W_A[2][27] = 4'hF;
    W_A[3][27] = 4'hF;
    W_A[4][27] = 4'hF;
    W_A[5][27] = 4'hF;
    W_A[6][27] = 4'hF;
    W_A[7][27] = 4'hF;
    W_A[8][27] = 4'hF;
    W_A[9][27] = 4'hF;
    W_A[10][27] = 4'hF;
    W_A[11][27] = 4'hF;
    W_A[12][27] = 4'hF;
    W_A[13][27] = 4'hF;
    W_A[14][27] = 4'hF;
    W_A[15][27] = 4'hF;
    W_A[16][27] = 4'hF;
    W_A[17][27] = 4'hF;
    W_A[18][27] = 4'hF;
    W_A[19][27] = 4'hF;
    W_A[20][27] = 4'hF;
    W_A[21][27] = 4'hF;
    W_A[22][27] = 4'hF;
    W_A[23][27] = 4'hF;
    W_A[24][27] = 4'hF;
    W_A[25][27] = 4'hF;
    W_A[26][27] = 4'hF;
    W_A[27][27] = 4'hF;
    W_A[28][27] = 4'hF;
    W_A[29][27] = 4'hF;
    W_A[30][27] = 4'hF;
    W_A[31][27] = 4'hF;
    W_A[32][27] = 4'hF;
    W_A[33][27] = 4'hF;
    W_A[34][27] = 4'hF;
    W_A[35][27] = 4'hF;
    W_A[36][27] = 4'hF;
    W_A[37][27] = 4'hF;
    W_A[38][27] = 4'hF;
    W_A[39][27] = 4'hF;
    W_A[40][27] = 4'hF;
    W_A[41][27] = 4'hF;
    W_A[42][27] = 4'hF;
    W_A[43][27] = 4'hF;
    W_A[44][27] = 4'hF;
    W_A[45][27] = 4'hF;
    W_A[46][27] = 4'hF;
    W_A[47][27] = 4'hF;
    W_A[48][27] = 4'hF;
    W_A[49][27] = 4'hF;
    W_A[50][27] = 4'hF;
    W_A[51][27] = 4'hF;
    W_A[52][27] = 4'hF;
    W_A[53][27] = 4'hF;
    W_A[54][27] = 4'hF;
    W_A[55][27] = 4'hF;
    W_A[56][27] = 4'hF;
    W_A[57][27] = 4'hF;
    W_A[58][27] = 4'hF;
    W_A[59][27] = 4'hF;
    W_A[60][27] = 4'hF;
    W_A[61][27] = 4'hF;
    W_A[62][27] = 4'hF;
    W_A[63][27] = 4'hF;
    W_A[64][27] = 4'hF;
    W_A[65][27] = 4'hF;
    W_A[66][27] = 4'hF;
    W_A[67][27] = 4'hF;
    W_A[68][27] = 4'hF;
    W_A[69][27] = 4'hF;
    W_A[70][27] = 4'hF;
    W_A[71][27] = 4'hF;
    W_A[72][27] = 4'hF;
    W_A[73][27] = 4'hF;
    W_A[74][27] = 4'hF;
    W_A[75][27] = 4'hF;
    W_A[76][27] = 4'hF;
    W_A[77][27] = 4'hF;
    W_A[78][27] = 4'hF;
    W_A[79][27] = 4'hF;
    W_A[80][27] = 4'hF;
    W_A[81][27] = 4'hF;
    W_A[82][27] = 4'hF;
    W_A[83][27] = 4'hF;
    W_A[84][27] = 4'hF;
    W_A[85][27] = 4'hF;
    W_A[86][27] = 4'hF;
    W_A[87][27] = 4'hF;
    W_A[88][27] = 4'hF;
    W_A[89][27] = 4'hF;
    W_A[90][27] = 4'hF;
    W_A[91][27] = 4'hF;
    W_A[92][27] = 4'hF;
    W_A[93][27] = 4'hF;
    W_A[94][27] = 4'hF;
    W_A[95][27] = 4'hF;
    W_A[96][27] = 4'hF;
    W_A[97][27] = 4'hF;
    W_A[98][27] = 4'hF;
    W_A[99][27] = 4'hF;
    W_A[100][27] = 4'hF;
    W_A[101][27] = 4'hF;
    W_A[102][27] = 4'hF;
    W_A[103][27] = 4'hF;
    W_A[104][27] = 4'hF;
    W_A[105][27] = 4'hF;
    W_A[106][27] = 4'hF;
    W_A[107][27] = 4'hF;
    W_A[0][28] = 4'hF;
    W_A[1][28] = 4'hF;
    W_A[2][28] = 4'hF;
    W_A[3][28] = 4'hF;
    W_A[4][28] = 4'hF;
    W_A[5][28] = 4'hF;
    W_A[6][28] = 4'hF;
    W_A[7][28] = 4'hF;
    W_A[8][28] = 4'hF;
    W_A[9][28] = 4'hF;
    W_A[10][28] = 4'hF;
    W_A[11][28] = 4'hF;
    W_A[12][28] = 4'hF;
    W_A[13][28] = 4'hF;
    W_A[14][28] = 4'hF;
    W_A[15][28] = 4'hF;
    W_A[16][28] = 4'hF;
    W_A[17][28] = 4'hF;
    W_A[18][28] = 4'hF;
    W_A[19][28] = 4'hF;
    W_A[20][28] = 4'hF;
    W_A[21][28] = 4'hF;
    W_A[22][28] = 4'hF;
    W_A[23][28] = 4'hF;
    W_A[24][28] = 4'hF;
    W_A[25][28] = 4'hF;
    W_A[26][28] = 4'hF;
    W_A[27][28] = 4'hF;
    W_A[28][28] = 4'hF;
    W_A[29][28] = 4'hF;
    W_A[30][28] = 4'hF;
    W_A[31][28] = 4'hF;
    W_A[32][28] = 4'hF;
    W_A[33][28] = 4'hF;
    W_A[34][28] = 4'hF;
    W_A[35][28] = 4'hF;
    W_A[36][28] = 4'hF;
    W_A[37][28] = 4'hF;
    W_A[38][28] = 4'hF;
    W_A[39][28] = 4'hF;
    W_A[40][28] = 4'hF;
    W_A[41][28] = 4'hF;
    W_A[42][28] = 4'hF;
    W_A[43][28] = 4'hF;
    W_A[44][28] = 4'hF;
    W_A[45][28] = 4'hF;
    W_A[46][28] = 4'hF;
    W_A[47][28] = 4'hF;
    W_A[48][28] = 4'hF;
    W_A[49][28] = 4'hF;
    W_A[50][28] = 4'hF;
    W_A[51][28] = 4'hF;
    W_A[52][28] = 4'hF;
    W_A[53][28] = 4'hF;
    W_A[54][28] = 4'hF;
    W_A[55][28] = 4'hF;
    W_A[56][28] = 4'hF;
    W_A[57][28] = 4'hF;
    W_A[58][28] = 4'hF;
    W_A[59][28] = 4'hF;
    W_A[60][28] = 4'hF;
    W_A[61][28] = 4'hF;
    W_A[62][28] = 4'hF;
    W_A[63][28] = 4'hF;
    W_A[64][28] = 4'hF;
    W_A[65][28] = 4'hF;
    W_A[66][28] = 4'hF;
    W_A[67][28] = 4'hF;
    W_A[68][28] = 4'hF;
    W_A[69][28] = 4'hF;
    W_A[70][28] = 4'hF;
    W_A[71][28] = 4'hF;
    W_A[72][28] = 4'hF;
    W_A[73][28] = 4'hF;
    W_A[74][28] = 4'hF;
    W_A[75][28] = 4'hF;
    W_A[76][28] = 4'hF;
    W_A[77][28] = 4'hF;
    W_A[78][28] = 4'hF;
    W_A[79][28] = 4'hF;
    W_A[80][28] = 4'hF;
    W_A[81][28] = 4'hF;
    W_A[82][28] = 4'hF;
    W_A[83][28] = 4'hF;
    W_A[84][28] = 4'hF;
    W_A[85][28] = 4'hF;
    W_A[86][28] = 4'hF;
    W_A[87][28] = 4'hF;
    W_A[88][28] = 4'hF;
    W_A[89][28] = 4'hF;
    W_A[90][28] = 4'hF;
    W_A[91][28] = 4'hF;
    W_A[92][28] = 4'hF;
    W_A[93][28] = 4'hF;
    W_A[94][28] = 4'hF;
    W_A[95][28] = 4'hF;
    W_A[96][28] = 4'hF;
    W_A[97][28] = 4'hF;
    W_A[98][28] = 4'hF;
    W_A[99][28] = 4'hF;
    W_A[100][28] = 4'hF;
    W_A[101][28] = 4'hF;
    W_A[102][28] = 4'hF;
    W_A[103][28] = 4'hF;
    W_A[104][28] = 4'hF;
    W_A[105][28] = 4'hF;
    W_A[106][28] = 4'hF;
    W_A[107][28] = 4'hF;

end

endmodule
