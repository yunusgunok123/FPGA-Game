module Numbers_init (
		output reg[3:0] Number0 [0:22][0:28],
		output reg[3:0] Number1 [0:22][0:28],
		output reg[3:0] Number2 [0:22][0:28],
		output reg[3:0] Number3 [0:22][0:28],
		output reg[3:0] Number4 [0:22][0:28],
		output reg[3:0] Number5 [0:22][0:28],
		output reg[3:0] Number6 [0:22][0:28],
		output reg[3:0] Number7 [0:22][0:28],
		output reg[3:0] Number8 [0:22][0:28],
		output reg[3:0] Number9 [0:22][0:28]

);
// Storing the pixel color information of Pictures of numbers for Score
initial begin
// Number 0
    Number0[0][0] = 4'hF;
    Number0[1][0] = 4'hF;
    Number0[2][0] = 4'hF;
    Number0[3][0] = 4'hF;
    Number0[4][0] = 4'hF;
    Number0[5][0] = 4'hF;
    Number0[6][0] = 4'hF;
    Number0[7][0] = 4'hF;
    Number0[8][0] = 4'hF;
    Number0[9][0] = 4'hF;
    Number0[10][0] = 4'hF;
    Number0[11][0] = 4'hF;
    Number0[12][0] = 4'hF;
    Number0[13][0] = 4'hF;
    Number0[14][0] = 4'hF;
    Number0[15][0] = 4'hF;
    Number0[16][0] = 4'hF;
    Number0[17][0] = 4'hF;
    Number0[18][0] = 4'hF;
    Number0[19][0] = 4'hF;
    Number0[20][0] = 4'hF;
    Number0[21][0] = 4'hF;
    Number0[22][0] = 4'hF;
    Number0[0][1] = 4'hF;
    Number0[1][1] = 4'hF;
    Number0[2][1] = 4'hF;
    Number0[3][1] = 4'hF;
    Number0[4][1] = 4'hF;
    Number0[5][1] = 4'hF;
    Number0[6][1] = 4'hF;
    Number0[7][1] = 4'hF;
    Number0[8][1] = 4'hF;
    Number0[9][1] = 4'hF;
    Number0[10][1] = 4'hF;
    Number0[11][1] = 4'hF;
    Number0[12][1] = 4'hF;
    Number0[13][1] = 4'hF;
    Number0[14][1] = 4'hF;
    Number0[15][1] = 4'hF;
    Number0[16][1] = 4'hF;
    Number0[17][1] = 4'hF;
    Number0[18][1] = 4'hF;
    Number0[19][1] = 4'hF;
    Number0[20][1] = 4'hF;
    Number0[21][1] = 4'hF;
    Number0[22][1] = 4'hF;
    Number0[0][2] = 4'hF;
    Number0[1][2] = 4'hF;
    Number0[2][2] = 4'hF;
    Number0[3][2] = 4'hF;
    Number0[4][2] = 4'hF;
    Number0[5][2] = 4'hF;
    Number0[6][2] = 4'hF;
    Number0[7][2] = 4'hE;
    Number0[8][2] = 4'hD;
    Number0[9][2] = 4'hC;
    Number0[10][2] = 4'hC;
    Number0[11][2] = 4'hC;
    Number0[12][2] = 4'hC;
    Number0[13][2] = 4'hC;
    Number0[14][2] = 4'hC;
    Number0[15][2] = 4'hD;
    Number0[16][2] = 4'hF;
    Number0[17][2] = 4'hF;
    Number0[18][2] = 4'hF;
    Number0[19][2] = 4'hF;
    Number0[20][2] = 4'hF;
    Number0[21][2] = 4'hF;
    Number0[22][2] = 4'hF;
    Number0[0][3] = 4'hF;
    Number0[1][3] = 4'hF;
    Number0[2][3] = 4'hF;
    Number0[3][3] = 4'hF;
    Number0[4][3] = 4'hF;
    Number0[5][3] = 4'hF;
    Number0[6][3] = 4'hD;
    Number0[7][3] = 4'hC;
    Number0[8][3] = 4'hC;
    Number0[9][3] = 4'hC;
    Number0[10][3] = 4'hC;
    Number0[11][3] = 4'hC;
    Number0[12][3] = 4'hC;
    Number0[13][3] = 4'hC;
    Number0[14][3] = 4'hC;
    Number0[15][3] = 4'hC;
    Number0[16][3] = 4'hC;
    Number0[17][3] = 4'hD;
    Number0[18][3] = 4'hF;
    Number0[19][3] = 4'hF;
    Number0[20][3] = 4'hF;
    Number0[21][3] = 4'hF;
    Number0[22][3] = 4'hF;
    Number0[0][4] = 4'hF;
    Number0[1][4] = 4'hF;
    Number0[2][4] = 4'hF;
    Number0[3][4] = 4'hF;
    Number0[4][4] = 4'hF;
    Number0[5][4] = 4'hD;
    Number0[6][4] = 4'hC;
    Number0[7][4] = 4'hC;
    Number0[8][4] = 4'hC;
    Number0[9][4] = 4'hC;
    Number0[10][4] = 4'hC;
    Number0[11][4] = 4'hC;
    Number0[12][4] = 4'hC;
    Number0[13][4] = 4'hC;
    Number0[14][4] = 4'hC;
    Number0[15][4] = 4'hC;
    Number0[16][4] = 4'hC;
    Number0[17][4] = 4'hC;
    Number0[18][4] = 4'hD;
    Number0[19][4] = 4'hF;
    Number0[20][4] = 4'hF;
    Number0[21][4] = 4'hF;
    Number0[22][4] = 4'hF;
    Number0[0][5] = 4'hF;
    Number0[1][5] = 4'hF;
    Number0[2][5] = 4'hF;
    Number0[3][5] = 4'hF;
    Number0[4][5] = 4'hD;
    Number0[5][5] = 4'hC;
    Number0[6][5] = 4'hC;
    Number0[7][5] = 4'hC;
    Number0[8][5] = 4'hC;
    Number0[9][5] = 4'hC;
    Number0[10][5] = 4'hC;
    Number0[11][5] = 4'hC;
    Number0[12][5] = 4'hC;
    Number0[13][5] = 4'hC;
    Number0[14][5] = 4'hC;
    Number0[15][5] = 4'hC;
    Number0[16][5] = 4'hC;
    Number0[17][5] = 4'hC;
    Number0[18][5] = 4'hC;
    Number0[19][5] = 4'hE;
    Number0[20][5] = 4'hF;
    Number0[21][5] = 4'hF;
    Number0[22][5] = 4'hF;
    Number0[0][6] = 4'hF;
    Number0[1][6] = 4'hF;
    Number0[2][6] = 4'hF;
    Number0[3][6] = 4'hF;
    Number0[4][6] = 4'hC;
    Number0[5][6] = 4'hC;
    Number0[6][6] = 4'hC;
    Number0[7][6] = 4'hC;
    Number0[8][6] = 4'hC;
    Number0[9][6] = 4'hC;
    Number0[10][6] = 4'hE;
    Number0[11][6] = 4'hF;
    Number0[12][6] = 4'hE;
    Number0[13][6] = 4'hD;
    Number0[14][6] = 4'hC;
    Number0[15][6] = 4'hC;
    Number0[16][6] = 4'hC;
    Number0[17][6] = 4'hC;
    Number0[18][6] = 4'hC;
    Number0[19][6] = 4'hD;
    Number0[20][6] = 4'hF;
    Number0[21][6] = 4'hF;
    Number0[22][6] = 4'hF;
    Number0[0][7] = 4'hF;
    Number0[1][7] = 4'hF;
    Number0[2][7] = 4'hF;
    Number0[3][7] = 4'hD;
    Number0[4][7] = 4'hC;
    Number0[5][7] = 4'hC;
    Number0[6][7] = 4'hC;
    Number0[7][7] = 4'hC;
    Number0[8][7] = 4'hC;
    Number0[9][7] = 4'hF;
    Number0[10][7] = 4'hF;
    Number0[11][7] = 4'hF;
    Number0[12][7] = 4'hF;
    Number0[13][7] = 4'hF;
    Number0[14][7] = 4'hD;
    Number0[15][7] = 4'hC;
    Number0[16][7] = 4'hC;
    Number0[17][7] = 4'hC;
    Number0[18][7] = 4'hC;
    Number0[19][7] = 4'hC;
    Number0[20][7] = 4'hF;
    Number0[21][7] = 4'hF;
    Number0[22][7] = 4'hF;
    Number0[0][8] = 4'hF;
    Number0[1][8] = 4'hF;
    Number0[2][8] = 4'hF;
    Number0[3][8] = 4'hD;
    Number0[4][8] = 4'hC;
    Number0[5][8] = 4'hC;
    Number0[6][8] = 4'hC;
    Number0[7][8] = 4'hC;
    Number0[8][8] = 4'hD;
    Number0[9][8] = 4'hF;
    Number0[10][8] = 4'hF;
    Number0[11][8] = 4'hF;
    Number0[12][8] = 4'hF;
    Number0[13][8] = 4'hF;
    Number0[14][8] = 4'hE;
    Number0[15][8] = 4'hC;
    Number0[16][8] = 4'hC;
    Number0[17][8] = 4'hC;
    Number0[18][8] = 4'hC;
    Number0[19][8] = 4'hC;
    Number0[20][8] = 4'hE;
    Number0[21][8] = 4'hF;
    Number0[22][8] = 4'hF;
    Number0[0][9] = 4'hF;
    Number0[1][9] = 4'hF;
    Number0[2][9] = 4'hF;
    Number0[3][9] = 4'hC;
    Number0[4][9] = 4'hC;
    Number0[5][9] = 4'hC;
    Number0[6][9] = 4'hC;
    Number0[7][9] = 4'hC;
    Number0[8][9] = 4'hE;
    Number0[9][9] = 4'hF;
    Number0[10][9] = 4'hF;
    Number0[11][9] = 4'hF;
    Number0[12][9] = 4'hF;
    Number0[13][9] = 4'hF;
    Number0[14][9] = 4'hF;
    Number0[15][9] = 4'hC;
    Number0[16][9] = 4'hC;
    Number0[17][9] = 4'hC;
    Number0[18][9] = 4'hC;
    Number0[19][9] = 4'hC;
    Number0[20][9] = 4'hD;
    Number0[21][9] = 4'hF;
    Number0[22][9] = 4'hF;
    Number0[0][10] = 4'hF;
    Number0[1][10] = 4'hF;
    Number0[2][10] = 4'hE;
    Number0[3][10] = 4'hC;
    Number0[4][10] = 4'hC;
    Number0[5][10] = 4'hC;
    Number0[6][10] = 4'hC;
    Number0[7][10] = 4'hC;
    Number0[8][10] = 4'hF;
    Number0[9][10] = 4'hF;
    Number0[10][10] = 4'hF;
    Number0[11][10] = 4'hF;
    Number0[12][10] = 4'hF;
    Number0[13][10] = 4'hF;
    Number0[14][10] = 4'hF;
    Number0[15][10] = 4'hC;
    Number0[16][10] = 4'hC;
    Number0[17][10] = 4'hC;
    Number0[18][10] = 4'hC;
    Number0[19][10] = 4'hC;
    Number0[20][10] = 4'hD;
    Number0[21][10] = 4'hF;
    Number0[22][10] = 4'hF;
    Number0[0][11] = 4'hF;
    Number0[1][11] = 4'hF;
    Number0[2][11] = 4'hE;
    Number0[3][11] = 4'hC;
    Number0[4][11] = 4'hC;
    Number0[5][11] = 4'hC;
    Number0[6][11] = 4'hC;
    Number0[7][11] = 4'hC;
    Number0[8][11] = 4'hF;
    Number0[9][11] = 4'hF;
    Number0[10][11] = 4'hF;
    Number0[11][11] = 4'hF;
    Number0[12][11] = 4'hF;
    Number0[13][11] = 4'hF;
    Number0[14][11] = 4'hF;
    Number0[15][11] = 4'hD;
    Number0[16][11] = 4'hC;
    Number0[17][11] = 4'hC;
    Number0[18][11] = 4'hC;
    Number0[19][11] = 4'hC;
    Number0[20][11] = 4'hD;
    Number0[21][11] = 4'hF;
    Number0[22][11] = 4'hF;
    Number0[0][12] = 4'hF;
    Number0[1][12] = 4'hF;
    Number0[2][12] = 4'hD;
    Number0[3][12] = 4'hC;
    Number0[4][12] = 4'hC;
    Number0[5][12] = 4'hC;
    Number0[6][12] = 4'hC;
    Number0[7][12] = 4'hC;
    Number0[8][12] = 4'hF;
    Number0[9][12] = 4'hF;
    Number0[10][12] = 4'hF;
    Number0[11][12] = 4'hF;
    Number0[12][12] = 4'hF;
    Number0[13][12] = 4'hF;
    Number0[14][12] = 4'hF;
    Number0[15][12] = 4'hD;
    Number0[16][12] = 4'hC;
    Number0[17][12] = 4'hC;
    Number0[18][12] = 4'hC;
    Number0[19][12] = 4'hC;
    Number0[20][12] = 4'hD;
    Number0[21][12] = 4'hF;
    Number0[22][12] = 4'hF;
    Number0[0][13] = 4'hF;
    Number0[1][13] = 4'hF;
    Number0[2][13] = 4'hD;
    Number0[3][13] = 4'hC;
    Number0[4][13] = 4'hC;
    Number0[5][13] = 4'hC;
    Number0[6][13] = 4'hC;
    Number0[7][13] = 4'hC;
    Number0[8][13] = 4'hF;
    Number0[9][13] = 4'hF;
    Number0[10][13] = 4'hF;
    Number0[11][13] = 4'hF;
    Number0[12][13] = 4'hF;
    Number0[13][13] = 4'hF;
    Number0[14][13] = 4'hF;
    Number0[15][13] = 4'hD;
    Number0[16][13] = 4'hC;
    Number0[17][13] = 4'hC;
    Number0[18][13] = 4'hC;
    Number0[19][13] = 4'hC;
    Number0[20][13] = 4'hD;
    Number0[21][13] = 4'hF;
    Number0[22][13] = 4'hF;
    Number0[0][14] = 4'hF;
    Number0[1][14] = 4'hF;
    Number0[2][14] = 4'hD;
    Number0[3][14] = 4'hC;
    Number0[4][14] = 4'hC;
    Number0[5][14] = 4'hC;
    Number0[6][14] = 4'hC;
    Number0[7][14] = 4'hC;
    Number0[8][14] = 4'hF;
    Number0[9][14] = 4'hF;
    Number0[10][14] = 4'hF;
    Number0[11][14] = 4'hF;
    Number0[12][14] = 4'hF;
    Number0[13][14] = 4'hF;
    Number0[14][14] = 4'hF;
    Number0[15][14] = 4'hD;
    Number0[16][14] = 4'hC;
    Number0[17][14] = 4'hC;
    Number0[18][14] = 4'hC;
    Number0[19][14] = 4'hC;
    Number0[20][14] = 4'hD;
    Number0[21][14] = 4'hF;
    Number0[22][14] = 4'hF;
    Number0[0][15] = 4'hF;
    Number0[1][15] = 4'hF;
    Number0[2][15] = 4'hD;
    Number0[3][15] = 4'hC;
    Number0[4][15] = 4'hC;
    Number0[5][15] = 4'hC;
    Number0[6][15] = 4'hC;
    Number0[7][15] = 4'hC;
    Number0[8][15] = 4'hF;
    Number0[9][15] = 4'hF;
    Number0[10][15] = 4'hF;
    Number0[11][15] = 4'hF;
    Number0[12][15] = 4'hF;
    Number0[13][15] = 4'hF;
    Number0[14][15] = 4'hF;
    Number0[15][15] = 4'hD;
    Number0[16][15] = 4'hC;
    Number0[17][15] = 4'hC;
    Number0[18][15] = 4'hC;
    Number0[19][15] = 4'hC;
    Number0[20][15] = 4'hD;
    Number0[21][15] = 4'hF;
    Number0[22][15] = 4'hF;
    Number0[0][16] = 4'hF;
    Number0[1][16] = 4'hF;
    Number0[2][16] = 4'hD;
    Number0[3][16] = 4'hC;
    Number0[4][16] = 4'hC;
    Number0[5][16] = 4'hC;
    Number0[6][16] = 4'hC;
    Number0[7][16] = 4'hC;
    Number0[8][16] = 4'hF;
    Number0[9][16] = 4'hF;
    Number0[10][16] = 4'hF;
    Number0[11][16] = 4'hF;
    Number0[12][16] = 4'hF;
    Number0[13][16] = 4'hF;
    Number0[14][16] = 4'hF;
    Number0[15][16] = 4'hD;
    Number0[16][16] = 4'hC;
    Number0[17][16] = 4'hC;
    Number0[18][16] = 4'hC;
    Number0[19][16] = 4'hC;
    Number0[20][16] = 4'hD;
    Number0[21][16] = 4'hF;
    Number0[22][16] = 4'hF;
    Number0[0][17] = 4'hF;
    Number0[1][17] = 4'hF;
    Number0[2][17] = 4'hD;
    Number0[3][17] = 4'hC;
    Number0[4][17] = 4'hC;
    Number0[5][17] = 4'hC;
    Number0[6][17] = 4'hC;
    Number0[7][17] = 4'hC;
    Number0[8][17] = 4'hF;
    Number0[9][17] = 4'hF;
    Number0[10][17] = 4'hF;
    Number0[11][17] = 4'hF;
    Number0[12][17] = 4'hF;
    Number0[13][17] = 4'hF;
    Number0[14][17] = 4'hF;
    Number0[15][17] = 4'hD;
    Number0[16][17] = 4'hC;
    Number0[17][17] = 4'hC;
    Number0[18][17] = 4'hC;
    Number0[19][17] = 4'hC;
    Number0[20][17] = 4'hD;
    Number0[21][17] = 4'hF;
    Number0[22][17] = 4'hF;
    Number0[0][18] = 4'hF;
    Number0[1][18] = 4'hF;
    Number0[2][18] = 4'hE;
    Number0[3][18] = 4'hC;
    Number0[4][18] = 4'hC;
    Number0[5][18] = 4'hC;
    Number0[6][18] = 4'hC;
    Number0[7][18] = 4'hC;
    Number0[8][18] = 4'hF;
    Number0[9][18] = 4'hF;
    Number0[10][18] = 4'hF;
    Number0[11][18] = 4'hF;
    Number0[12][18] = 4'hF;
    Number0[13][18] = 4'hF;
    Number0[14][18] = 4'hF;
    Number0[15][18] = 4'hC;
    Number0[16][18] = 4'hC;
    Number0[17][18] = 4'hC;
    Number0[18][18] = 4'hC;
    Number0[19][18] = 4'hC;
    Number0[20][18] = 4'hD;
    Number0[21][18] = 4'hF;
    Number0[22][18] = 4'hF;
    Number0[0][19] = 4'hF;
    Number0[1][19] = 4'hF;
    Number0[2][19] = 4'hF;
    Number0[3][19] = 4'hC;
    Number0[4][19] = 4'hC;
    Number0[5][19] = 4'hC;
    Number0[6][19] = 4'hC;
    Number0[7][19] = 4'hC;
    Number0[8][19] = 4'hE;
    Number0[9][19] = 4'hF;
    Number0[10][19] = 4'hF;
    Number0[11][19] = 4'hF;
    Number0[12][19] = 4'hF;
    Number0[13][19] = 4'hF;
    Number0[14][19] = 4'hF;
    Number0[15][19] = 4'hC;
    Number0[16][19] = 4'hC;
    Number0[17][19] = 4'hC;
    Number0[18][19] = 4'hC;
    Number0[19][19] = 4'hC;
    Number0[20][19] = 4'hE;
    Number0[21][19] = 4'hF;
    Number0[22][19] = 4'hF;
    Number0[0][20] = 4'hF;
    Number0[1][20] = 4'hF;
    Number0[2][20] = 4'hF;
    Number0[3][20] = 4'hC;
    Number0[4][20] = 4'hC;
    Number0[5][20] = 4'hC;
    Number0[6][20] = 4'hC;
    Number0[7][20] = 4'hC;
    Number0[8][20] = 4'hD;
    Number0[9][20] = 4'hF;
    Number0[10][20] = 4'hF;
    Number0[11][20] = 4'hF;
    Number0[12][20] = 4'hF;
    Number0[13][20] = 4'hF;
    Number0[14][20] = 4'hE;
    Number0[15][20] = 4'hC;
    Number0[16][20] = 4'hC;
    Number0[17][20] = 4'hC;
    Number0[18][20] = 4'hC;
    Number0[19][20] = 4'hC;
    Number0[20][20] = 4'hF;
    Number0[21][20] = 4'hF;
    Number0[22][20] = 4'hF;
    Number0[0][21] = 4'hF;
    Number0[1][21] = 4'hF;
    Number0[2][21] = 4'hF;
    Number0[3][21] = 4'hD;
    Number0[4][21] = 4'hC;
    Number0[5][21] = 4'hC;
    Number0[6][21] = 4'hC;
    Number0[7][21] = 4'hC;
    Number0[8][21] = 4'hC;
    Number0[9][21] = 4'hF;
    Number0[10][21] = 4'hF;
    Number0[11][21] = 4'hF;
    Number0[12][21] = 4'hF;
    Number0[13][21] = 4'hF;
    Number0[14][21] = 4'hD;
    Number0[15][21] = 4'hC;
    Number0[16][21] = 4'hC;
    Number0[17][21] = 4'hC;
    Number0[18][21] = 4'hC;
    Number0[19][21] = 4'hD;
    Number0[20][21] = 4'hF;
    Number0[21][21] = 4'hF;
    Number0[22][21] = 4'hF;
    Number0[0][22] = 4'hF;
    Number0[1][22] = 4'hF;
    Number0[2][22] = 4'hF;
    Number0[3][22] = 4'hE;
    Number0[4][22] = 4'hC;
    Number0[5][22] = 4'hC;
    Number0[6][22] = 4'hC;
    Number0[7][22] = 4'hC;
    Number0[8][22] = 4'hC;
    Number0[9][22] = 4'hD;
    Number0[10][22] = 4'hE;
    Number0[11][22] = 4'hF;
    Number0[12][22] = 4'hE;
    Number0[13][22] = 4'hD;
    Number0[14][22] = 4'hC;
    Number0[15][22] = 4'hC;
    Number0[16][22] = 4'hC;
    Number0[17][22] = 4'hC;
    Number0[18][22] = 4'hC;
    Number0[19][22] = 4'hE;
    Number0[20][22] = 4'hF;
    Number0[21][22] = 4'hF;
    Number0[22][22] = 4'hF;
    Number0[0][23] = 4'hF;
    Number0[1][23] = 4'hF;
    Number0[2][23] = 4'hF;
    Number0[3][23] = 4'hF;
    Number0[4][23] = 4'hD;
    Number0[5][23] = 4'hC;
    Number0[6][23] = 4'hC;
    Number0[7][23] = 4'hC;
    Number0[8][23] = 4'hC;
    Number0[9][23] = 4'hC;
    Number0[10][23] = 4'hC;
    Number0[11][23] = 4'hC;
    Number0[12][23] = 4'hC;
    Number0[13][23] = 4'hC;
    Number0[14][23] = 4'hC;
    Number0[15][23] = 4'hC;
    Number0[16][23] = 4'hC;
    Number0[17][23] = 4'hC;
    Number0[18][23] = 4'hD;
    Number0[19][23] = 4'hF;
    Number0[20][23] = 4'hF;
    Number0[21][23] = 4'hF;
    Number0[22][23] = 4'hF;
    Number0[0][24] = 4'hF;
    Number0[1][24] = 4'hF;
    Number0[2][24] = 4'hF;
    Number0[3][24] = 4'hF;
    Number0[4][24] = 4'hE;
    Number0[5][24] = 4'hC;
    Number0[6][24] = 4'hC;
    Number0[7][24] = 4'hC;
    Number0[8][24] = 4'hC;
    Number0[9][24] = 4'hC;
    Number0[10][24] = 4'hC;
    Number0[11][24] = 4'hC;
    Number0[12][24] = 4'hC;
    Number0[13][24] = 4'hC;
    Number0[14][24] = 4'hC;
    Number0[15][24] = 4'hC;
    Number0[16][24] = 4'hC;
    Number0[17][24] = 4'hC;
    Number0[18][24] = 4'hF;
    Number0[19][24] = 4'hF;
    Number0[20][24] = 4'hF;
    Number0[21][24] = 4'hF;
    Number0[22][24] = 4'hF;
    Number0[0][25] = 4'hF;
    Number0[1][25] = 4'hF;
    Number0[2][25] = 4'hF;
    Number0[3][25] = 4'hF;
    Number0[4][25] = 4'hF;
    Number0[5][25] = 4'hE;
    Number0[6][25] = 4'hC;
    Number0[7][25] = 4'hC;
    Number0[8][25] = 4'hC;
    Number0[9][25] = 4'hC;
    Number0[10][25] = 4'hC;
    Number0[11][25] = 4'hC;
    Number0[12][25] = 4'hC;
    Number0[13][25] = 4'hC;
    Number0[14][25] = 4'hC;
    Number0[15][25] = 4'hC;
    Number0[16][25] = 4'hD;
    Number0[17][25] = 4'hE;
    Number0[18][25] = 4'hF;
    Number0[19][25] = 4'hF;
    Number0[20][25] = 4'hF;
    Number0[21][25] = 4'hF;
    Number0[22][25] = 4'hF;
    Number0[0][26] = 4'hF;
    Number0[1][26] = 4'hF;
    Number0[2][26] = 4'hF;
    Number0[3][26] = 4'hF;
    Number0[4][26] = 4'hF;
    Number0[5][26] = 4'hF;
    Number0[6][26] = 4'hF;
    Number0[7][26] = 4'hD;
    Number0[8][26] = 4'hD;
    Number0[9][26] = 4'hC;
    Number0[10][26] = 4'hC;
    Number0[11][26] = 4'hC;
    Number0[12][26] = 4'hC;
    Number0[13][26] = 4'hC;
    Number0[14][26] = 4'hD;
    Number0[15][26] = 4'hE;
    Number0[16][26] = 4'hF;
    Number0[17][26] = 4'hF;
    Number0[18][26] = 4'hF;
    Number0[19][26] = 4'hF;
    Number0[20][26] = 4'hF;
    Number0[21][26] = 4'hF;
    Number0[22][26] = 4'hF;
    Number0[0][27] = 4'hF;
    Number0[1][27] = 4'hF;
    Number0[2][27] = 4'hF;
    Number0[3][27] = 4'hF;
    Number0[4][27] = 4'hF;
    Number0[5][27] = 4'hF;
    Number0[6][27] = 4'hF;
    Number0[7][27] = 4'hF;
    Number0[8][27] = 4'hF;
    Number0[9][27] = 4'hF;
    Number0[10][27] = 4'hF;
    Number0[11][27] = 4'hF;
    Number0[12][27] = 4'hF;
    Number0[13][27] = 4'hF;
    Number0[14][27] = 4'hF;
    Number0[15][27] = 4'hF;
    Number0[16][27] = 4'hF;
    Number0[17][27] = 4'hF;
    Number0[18][27] = 4'hF;
    Number0[19][27] = 4'hF;
    Number0[20][27] = 4'hF;
    Number0[21][27] = 4'hF;
    Number0[22][27] = 4'hF;
    Number0[0][28] = 4'hF;
    Number0[1][28] = 4'hF;
    Number0[2][28] = 4'hF;
    Number0[3][28] = 4'hF;
    Number0[4][28] = 4'hF;
    Number0[5][28] = 4'hF;
    Number0[6][28] = 4'hF;
    Number0[7][28] = 4'hF;
    Number0[8][28] = 4'hF;
    Number0[9][28] = 4'hF;
    Number0[10][28] = 4'hF;
    Number0[11][28] = 4'hF;
    Number0[12][28] = 4'hF;
    Number0[13][28] = 4'hF;
    Number0[14][28] = 4'hF;
    Number0[15][28] = 4'hF;
    Number0[16][28] = 4'hF;
    Number0[17][28] = 4'hF;
    Number0[18][28] = 4'hF;
    Number0[19][28] = 4'hF;
    Number0[20][28] = 4'hF;
    Number0[21][28] = 4'hF;
    Number0[22][28] = 4'hF;

// Number 1
    Number1[0][0] = 4'hF;
    Number1[1][0] = 4'hF;
    Number1[2][0] = 4'hF;
    Number1[3][0] = 4'hF;
    Number1[4][0] = 4'hF;
    Number1[5][0] = 4'hF;
    Number1[6][0] = 4'hF;
    Number1[7][0] = 4'hF;
    Number1[8][0] = 4'hF;
    Number1[9][0] = 4'hF;
    Number1[10][0] = 4'hF;
    Number1[11][0] = 4'hF;
    Number1[12][0] = 4'hF;
    Number1[13][0] = 4'hF;
    Number1[14][0] = 4'hF;
    Number1[15][0] = 4'hF;
    Number1[16][0] = 4'hF;
    Number1[17][0] = 4'hF;
    Number1[18][0] = 4'hF;
    Number1[19][0] = 4'hF;
    Number1[20][0] = 4'hF;
    Number1[21][0] = 4'hF;
    Number1[22][0] = 4'hF;
    Number1[0][1] = 4'hF;
    Number1[1][1] = 4'hF;
    Number1[2][1] = 4'hF;
    Number1[3][1] = 4'hF;
    Number1[4][1] = 4'hF;
    Number1[5][1] = 4'hF;
    Number1[6][1] = 4'hF;
    Number1[7][1] = 4'hF;
    Number1[8][1] = 4'hF;
    Number1[9][1] = 4'hF;
    Number1[10][1] = 4'hF;
    Number1[11][1] = 4'hF;
    Number1[12][1] = 4'hF;
    Number1[13][1] = 4'hF;
    Number1[14][1] = 4'hF;
    Number1[15][1] = 4'hF;
    Number1[16][1] = 4'hF;
    Number1[17][1] = 4'hF;
    Number1[18][1] = 4'hF;
    Number1[19][1] = 4'hF;
    Number1[20][1] = 4'hF;
    Number1[21][1] = 4'hF;
    Number1[22][1] = 4'hF;
    Number1[0][2] = 4'hF;
    Number1[1][2] = 4'hF;
    Number1[2][2] = 4'hF;
    Number1[3][2] = 4'hF;
    Number1[4][2] = 4'hF;
    Number1[5][2] = 4'hF;
    Number1[6][2] = 4'hF;
    Number1[7][2] = 4'hF;
    Number1[8][2] = 4'hF;
    Number1[9][2] = 4'hE;
    Number1[10][2] = 4'hC;
    Number1[11][2] = 4'hC;
    Number1[12][2] = 4'hC;
    Number1[13][2] = 4'hC;
    Number1[14][2] = 4'hC;
    Number1[15][2] = 4'hF;
    Number1[16][2] = 4'hF;
    Number1[17][2] = 4'hF;
    Number1[18][2] = 4'hF;
    Number1[19][2] = 4'hF;
    Number1[20][2] = 4'hF;
    Number1[21][2] = 4'hF;
    Number1[22][2] = 4'hF;
    Number1[0][3] = 4'hF;
    Number1[1][3] = 4'hF;
    Number1[2][3] = 4'hF;
    Number1[3][3] = 4'hF;
    Number1[4][3] = 4'hF;
    Number1[5][3] = 4'hF;
    Number1[6][3] = 4'hF;
    Number1[7][3] = 4'hF;
    Number1[8][3] = 4'hD;
    Number1[9][3] = 4'hC;
    Number1[10][3] = 4'hC;
    Number1[11][3] = 4'hC;
    Number1[12][3] = 4'hC;
    Number1[13][3] = 4'hC;
    Number1[14][3] = 4'hC;
    Number1[15][3] = 4'hF;
    Number1[16][3] = 4'hF;
    Number1[17][3] = 4'hF;
    Number1[18][3] = 4'hF;
    Number1[19][3] = 4'hF;
    Number1[20][3] = 4'hF;
    Number1[21][3] = 4'hF;
    Number1[22][3] = 4'hF;
    Number1[0][4] = 4'hF;
    Number1[1][4] = 4'hF;
    Number1[2][4] = 4'hF;
    Number1[3][4] = 4'hF;
    Number1[4][4] = 4'hF;
    Number1[5][4] = 4'hF;
    Number1[6][4] = 4'hD;
    Number1[7][4] = 4'hC;
    Number1[8][4] = 4'hC;
    Number1[9][4] = 4'hC;
    Number1[10][4] = 4'hC;
    Number1[11][4] = 4'hC;
    Number1[12][4] = 4'hC;
    Number1[13][4] = 4'hC;
    Number1[14][4] = 4'hC;
    Number1[15][4] = 4'hF;
    Number1[16][4] = 4'hF;
    Number1[17][4] = 4'hF;
    Number1[18][4] = 4'hF;
    Number1[19][4] = 4'hF;
    Number1[20][4] = 4'hF;
    Number1[21][4] = 4'hF;
    Number1[22][4] = 4'hF;
    Number1[0][5] = 4'hF;
    Number1[1][5] = 4'hF;
    Number1[2][5] = 4'hF;
    Number1[3][5] = 4'hF;
    Number1[4][5] = 4'hE;
    Number1[5][5] = 4'hD;
    Number1[6][5] = 4'hC;
    Number1[7][5] = 4'hC;
    Number1[8][5] = 4'hC;
    Number1[9][5] = 4'hC;
    Number1[10][5] = 4'hC;
    Number1[11][5] = 4'hC;
    Number1[12][5] = 4'hC;
    Number1[13][5] = 4'hC;
    Number1[14][5] = 4'hC;
    Number1[15][5] = 4'hF;
    Number1[16][5] = 4'hF;
    Number1[17][5] = 4'hF;
    Number1[18][5] = 4'hF;
    Number1[19][5] = 4'hF;
    Number1[20][5] = 4'hF;
    Number1[21][5] = 4'hF;
    Number1[22][5] = 4'hF;
    Number1[0][6] = 4'hF;
    Number1[1][6] = 4'hF;
    Number1[2][6] = 4'hF;
    Number1[3][6] = 4'hF;
    Number1[4][6] = 4'hD;
    Number1[5][6] = 4'hC;
    Number1[6][6] = 4'hC;
    Number1[7][6] = 4'hC;
    Number1[8][6] = 4'hC;
    Number1[9][6] = 4'hC;
    Number1[10][6] = 4'hC;
    Number1[11][6] = 4'hC;
    Number1[12][6] = 4'hC;
    Number1[13][6] = 4'hC;
    Number1[14][6] = 4'hC;
    Number1[15][6] = 4'hF;
    Number1[16][6] = 4'hF;
    Number1[17][6] = 4'hF;
    Number1[18][6] = 4'hF;
    Number1[19][6] = 4'hF;
    Number1[20][6] = 4'hF;
    Number1[21][6] = 4'hF;
    Number1[22][6] = 4'hF;
    Number1[0][7] = 4'hF;
    Number1[1][7] = 4'hF;
    Number1[2][7] = 4'hF;
    Number1[3][7] = 4'hF;
    Number1[4][7] = 4'hD;
    Number1[5][7] = 4'hC;
    Number1[6][7] = 4'hC;
    Number1[7][7] = 4'hC;
    Number1[8][7] = 4'hC;
    Number1[9][7] = 4'hD;
    Number1[10][7] = 4'hC;
    Number1[11][7] = 4'hC;
    Number1[12][7] = 4'hC;
    Number1[13][7] = 4'hC;
    Number1[14][7] = 4'hC;
    Number1[15][7] = 4'hF;
    Number1[16][7] = 4'hF;
    Number1[17][7] = 4'hF;
    Number1[18][7] = 4'hF;
    Number1[19][7] = 4'hF;
    Number1[20][7] = 4'hF;
    Number1[21][7] = 4'hF;
    Number1[22][7] = 4'hF;
    Number1[0][8] = 4'hF;
    Number1[1][8] = 4'hF;
    Number1[2][8] = 4'hF;
    Number1[3][8] = 4'hF;
    Number1[4][8] = 4'hD;
    Number1[5][8] = 4'hC;
    Number1[6][8] = 4'hD;
    Number1[7][8] = 4'hE;
    Number1[8][8] = 4'hF;
    Number1[9][8] = 4'hE;
    Number1[10][8] = 4'hC;
    Number1[11][8] = 4'hC;
    Number1[12][8] = 4'hC;
    Number1[13][8] = 4'hC;
    Number1[14][8] = 4'hC;
    Number1[15][8] = 4'hF;
    Number1[16][8] = 4'hF;
    Number1[17][8] = 4'hF;
    Number1[18][8] = 4'hF;
    Number1[19][8] = 4'hF;
    Number1[20][8] = 4'hF;
    Number1[21][8] = 4'hF;
    Number1[22][8] = 4'hF;
    Number1[0][9] = 4'hF;
    Number1[1][9] = 4'hF;
    Number1[2][9] = 4'hF;
    Number1[3][9] = 4'hF;
    Number1[4][9] = 4'hE;
    Number1[5][9] = 4'hE;
    Number1[6][9] = 4'hF;
    Number1[7][9] = 4'hF;
    Number1[8][9] = 4'hF;
    Number1[9][9] = 4'hE;
    Number1[10][9] = 4'hC;
    Number1[11][9] = 4'hC;
    Number1[12][9] = 4'hC;
    Number1[13][9] = 4'hC;
    Number1[14][9] = 4'hC;
    Number1[15][9] = 4'hF;
    Number1[16][9] = 4'hF;
    Number1[17][9] = 4'hF;
    Number1[18][9] = 4'hF;
    Number1[19][9] = 4'hF;
    Number1[20][9] = 4'hF;
    Number1[21][9] = 4'hF;
    Number1[22][9] = 4'hF;
    Number1[0][10] = 4'hF;
    Number1[1][10] = 4'hF;
    Number1[2][10] = 4'hF;
    Number1[3][10] = 4'hF;
    Number1[4][10] = 4'hF;
    Number1[5][10] = 4'hF;
    Number1[6][10] = 4'hF;
    Number1[7][10] = 4'hF;
    Number1[8][10] = 4'hF;
    Number1[9][10] = 4'hE;
    Number1[10][10] = 4'hC;
    Number1[11][10] = 4'hC;
    Number1[12][10] = 4'hC;
    Number1[13][10] = 4'hC;
    Number1[14][10] = 4'hC;
    Number1[15][10] = 4'hF;
    Number1[16][10] = 4'hF;
    Number1[17][10] = 4'hF;
    Number1[18][10] = 4'hF;
    Number1[19][10] = 4'hF;
    Number1[20][10] = 4'hF;
    Number1[21][10] = 4'hF;
    Number1[22][10] = 4'hF;
    Number1[0][11] = 4'hF;
    Number1[1][11] = 4'hF;
    Number1[2][11] = 4'hF;
    Number1[3][11] = 4'hF;
    Number1[4][11] = 4'hF;
    Number1[5][11] = 4'hF;
    Number1[6][11] = 4'hF;
    Number1[7][11] = 4'hF;
    Number1[8][11] = 4'hF;
    Number1[9][11] = 4'hE;
    Number1[10][11] = 4'hC;
    Number1[11][11] = 4'hC;
    Number1[12][11] = 4'hC;
    Number1[13][11] = 4'hC;
    Number1[14][11] = 4'hC;
    Number1[15][11] = 4'hF;
    Number1[16][11] = 4'hF;
    Number1[17][11] = 4'hF;
    Number1[18][11] = 4'hF;
    Number1[19][11] = 4'hF;
    Number1[20][11] = 4'hF;
    Number1[21][11] = 4'hF;
    Number1[22][11] = 4'hF;
    Number1[0][12] = 4'hF;
    Number1[1][12] = 4'hF;
    Number1[2][12] = 4'hF;
    Number1[3][12] = 4'hF;
    Number1[4][12] = 4'hF;
    Number1[5][12] = 4'hF;
    Number1[6][12] = 4'hF;
    Number1[7][12] = 4'hF;
    Number1[8][12] = 4'hF;
    Number1[9][12] = 4'hE;
    Number1[10][12] = 4'hC;
    Number1[11][12] = 4'hC;
    Number1[12][12] = 4'hC;
    Number1[13][12] = 4'hC;
    Number1[14][12] = 4'hC;
    Number1[15][12] = 4'hF;
    Number1[16][12] = 4'hF;
    Number1[17][12] = 4'hF;
    Number1[18][12] = 4'hF;
    Number1[19][12] = 4'hF;
    Number1[20][12] = 4'hF;
    Number1[21][12] = 4'hF;
    Number1[22][12] = 4'hF;
    Number1[0][13] = 4'hF;
    Number1[1][13] = 4'hF;
    Number1[2][13] = 4'hF;
    Number1[3][13] = 4'hF;
    Number1[4][13] = 4'hF;
    Number1[5][13] = 4'hF;
    Number1[6][13] = 4'hF;
    Number1[7][13] = 4'hF;
    Number1[8][13] = 4'hF;
    Number1[9][13] = 4'hE;
    Number1[10][13] = 4'hC;
    Number1[11][13] = 4'hC;
    Number1[12][13] = 4'hC;
    Number1[13][13] = 4'hC;
    Number1[14][13] = 4'hC;
    Number1[15][13] = 4'hF;
    Number1[16][13] = 4'hF;
    Number1[17][13] = 4'hF;
    Number1[18][13] = 4'hF;
    Number1[19][13] = 4'hF;
    Number1[20][13] = 4'hF;
    Number1[21][13] = 4'hF;
    Number1[22][13] = 4'hF;
    Number1[0][14] = 4'hF;
    Number1[1][14] = 4'hF;
    Number1[2][14] = 4'hF;
    Number1[3][14] = 4'hF;
    Number1[4][14] = 4'hF;
    Number1[5][14] = 4'hF;
    Number1[6][14] = 4'hF;
    Number1[7][14] = 4'hF;
    Number1[8][14] = 4'hF;
    Number1[9][14] = 4'hE;
    Number1[10][14] = 4'hC;
    Number1[11][14] = 4'hC;
    Number1[12][14] = 4'hC;
    Number1[13][14] = 4'hC;
    Number1[14][14] = 4'hC;
    Number1[15][14] = 4'hF;
    Number1[16][14] = 4'hF;
    Number1[17][14] = 4'hF;
    Number1[18][14] = 4'hF;
    Number1[19][14] = 4'hF;
    Number1[20][14] = 4'hF;
    Number1[21][14] = 4'hF;
    Number1[22][14] = 4'hF;
    Number1[0][15] = 4'hF;
    Number1[1][15] = 4'hF;
    Number1[2][15] = 4'hF;
    Number1[3][15] = 4'hF;
    Number1[4][15] = 4'hF;
    Number1[5][15] = 4'hF;
    Number1[6][15] = 4'hF;
    Number1[7][15] = 4'hF;
    Number1[8][15] = 4'hF;
    Number1[9][15] = 4'hE;
    Number1[10][15] = 4'hC;
    Number1[11][15] = 4'hC;
    Number1[12][15] = 4'hC;
    Number1[13][15] = 4'hC;
    Number1[14][15] = 4'hC;
    Number1[15][15] = 4'hF;
    Number1[16][15] = 4'hF;
    Number1[17][15] = 4'hF;
    Number1[18][15] = 4'hF;
    Number1[19][15] = 4'hF;
    Number1[20][15] = 4'hF;
    Number1[21][15] = 4'hF;
    Number1[22][15] = 4'hF;
    Number1[0][16] = 4'hF;
    Number1[1][16] = 4'hF;
    Number1[2][16] = 4'hF;
    Number1[3][16] = 4'hF;
    Number1[4][16] = 4'hF;
    Number1[5][16] = 4'hF;
    Number1[6][16] = 4'hF;
    Number1[7][16] = 4'hF;
    Number1[8][16] = 4'hF;
    Number1[9][16] = 4'hE;
    Number1[10][16] = 4'hC;
    Number1[11][16] = 4'hC;
    Number1[12][16] = 4'hC;
    Number1[13][16] = 4'hC;
    Number1[14][16] = 4'hC;
    Number1[15][16] = 4'hF;
    Number1[16][16] = 4'hF;
    Number1[17][16] = 4'hF;
    Number1[18][16] = 4'hF;
    Number1[19][16] = 4'hF;
    Number1[20][16] = 4'hF;
    Number1[21][16] = 4'hF;
    Number1[22][16] = 4'hF;
    Number1[0][17] = 4'hF;
    Number1[1][17] = 4'hF;
    Number1[2][17] = 4'hF;
    Number1[3][17] = 4'hF;
    Number1[4][17] = 4'hF;
    Number1[5][17] = 4'hF;
    Number1[6][17] = 4'hF;
    Number1[7][17] = 4'hF;
    Number1[8][17] = 4'hF;
    Number1[9][17] = 4'hE;
    Number1[10][17] = 4'hC;
    Number1[11][17] = 4'hC;
    Number1[12][17] = 4'hC;
    Number1[13][17] = 4'hC;
    Number1[14][17] = 4'hC;
    Number1[15][17] = 4'hF;
    Number1[16][17] = 4'hF;
    Number1[17][17] = 4'hF;
    Number1[18][17] = 4'hF;
    Number1[19][17] = 4'hF;
    Number1[20][17] = 4'hF;
    Number1[21][17] = 4'hF;
    Number1[22][17] = 4'hF;
    Number1[0][18] = 4'hF;
    Number1[1][18] = 4'hF;
    Number1[2][18] = 4'hF;
    Number1[3][18] = 4'hF;
    Number1[4][18] = 4'hF;
    Number1[5][18] = 4'hF;
    Number1[6][18] = 4'hF;
    Number1[7][18] = 4'hF;
    Number1[8][18] = 4'hF;
    Number1[9][18] = 4'hE;
    Number1[10][18] = 4'hC;
    Number1[11][18] = 4'hC;
    Number1[12][18] = 4'hC;
    Number1[13][18] = 4'hC;
    Number1[14][18] = 4'hC;
    Number1[15][18] = 4'hF;
    Number1[16][18] = 4'hF;
    Number1[17][18] = 4'hF;
    Number1[18][18] = 4'hF;
    Number1[19][18] = 4'hF;
    Number1[20][18] = 4'hF;
    Number1[21][18] = 4'hF;
    Number1[22][18] = 4'hF;
    Number1[0][19] = 4'hF;
    Number1[1][19] = 4'hF;
    Number1[2][19] = 4'hF;
    Number1[3][19] = 4'hF;
    Number1[4][19] = 4'hF;
    Number1[5][19] = 4'hF;
    Number1[6][19] = 4'hF;
    Number1[7][19] = 4'hF;
    Number1[8][19] = 4'hF;
    Number1[9][19] = 4'hE;
    Number1[10][19] = 4'hC;
    Number1[11][19] = 4'hC;
    Number1[12][19] = 4'hC;
    Number1[13][19] = 4'hC;
    Number1[14][19] = 4'hC;
    Number1[15][19] = 4'hF;
    Number1[16][19] = 4'hF;
    Number1[17][19] = 4'hF;
    Number1[18][19] = 4'hF;
    Number1[19][19] = 4'hF;
    Number1[20][19] = 4'hF;
    Number1[21][19] = 4'hF;
    Number1[22][19] = 4'hF;
    Number1[0][20] = 4'hF;
    Number1[1][20] = 4'hF;
    Number1[2][20] = 4'hF;
    Number1[3][20] = 4'hF;
    Number1[4][20] = 4'hF;
    Number1[5][20] = 4'hF;
    Number1[6][20] = 4'hF;
    Number1[7][20] = 4'hF;
    Number1[8][20] = 4'hF;
    Number1[9][20] = 4'hE;
    Number1[10][20] = 4'hC;
    Number1[11][20] = 4'hC;
    Number1[12][20] = 4'hC;
    Number1[13][20] = 4'hC;
    Number1[14][20] = 4'hC;
    Number1[15][20] = 4'hF;
    Number1[16][20] = 4'hF;
    Number1[17][20] = 4'hF;
    Number1[18][20] = 4'hF;
    Number1[19][20] = 4'hF;
    Number1[20][20] = 4'hF;
    Number1[21][20] = 4'hF;
    Number1[22][20] = 4'hF;
    Number1[0][21] = 4'hF;
    Number1[1][21] = 4'hF;
    Number1[2][21] = 4'hF;
    Number1[3][21] = 4'hF;
    Number1[4][21] = 4'hF;
    Number1[5][21] = 4'hF;
    Number1[6][21] = 4'hF;
    Number1[7][21] = 4'hF;
    Number1[8][21] = 4'hF;
    Number1[9][21] = 4'hE;
    Number1[10][21] = 4'hC;
    Number1[11][21] = 4'hC;
    Number1[12][21] = 4'hC;
    Number1[13][21] = 4'hC;
    Number1[14][21] = 4'hC;
    Number1[15][21] = 4'hF;
    Number1[16][21] = 4'hF;
    Number1[17][21] = 4'hF;
    Number1[18][21] = 4'hF;
    Number1[19][21] = 4'hF;
    Number1[20][21] = 4'hF;
    Number1[21][21] = 4'hF;
    Number1[22][21] = 4'hF;
    Number1[0][22] = 4'hF;
    Number1[1][22] = 4'hF;
    Number1[2][22] = 4'hF;
    Number1[3][22] = 4'hF;
    Number1[4][22] = 4'hF;
    Number1[5][22] = 4'hF;
    Number1[6][22] = 4'hF;
    Number1[7][22] = 4'hF;
    Number1[8][22] = 4'hF;
    Number1[9][22] = 4'hE;
    Number1[10][22] = 4'hC;
    Number1[11][22] = 4'hC;
    Number1[12][22] = 4'hC;
    Number1[13][22] = 4'hC;
    Number1[14][22] = 4'hC;
    Number1[15][22] = 4'hF;
    Number1[16][22] = 4'hF;
    Number1[17][22] = 4'hF;
    Number1[18][22] = 4'hF;
    Number1[19][22] = 4'hF;
    Number1[20][22] = 4'hF;
    Number1[21][22] = 4'hF;
    Number1[22][22] = 4'hF;
    Number1[0][23] = 4'hF;
    Number1[1][23] = 4'hF;
    Number1[2][23] = 4'hF;
    Number1[3][23] = 4'hF;
    Number1[4][23] = 4'hD;
    Number1[5][23] = 4'hC;
    Number1[6][23] = 4'hC;
    Number1[7][23] = 4'hC;
    Number1[8][23] = 4'hC;
    Number1[9][23] = 4'hC;
    Number1[10][23] = 4'hC;
    Number1[11][23] = 4'hC;
    Number1[12][23] = 4'hC;
    Number1[13][23] = 4'hC;
    Number1[14][23] = 4'hC;
    Number1[15][23] = 4'hC;
    Number1[16][23] = 4'hC;
    Number1[17][23] = 4'hC;
    Number1[18][23] = 4'hC;
    Number1[19][23] = 4'hD;
    Number1[20][23] = 4'hF;
    Number1[21][23] = 4'hF;
    Number1[22][23] = 4'hF;
    Number1[0][24] = 4'hF;
    Number1[1][24] = 4'hF;
    Number1[2][24] = 4'hF;
    Number1[3][24] = 4'hF;
    Number1[4][24] = 4'hD;
    Number1[5][24] = 4'hC;
    Number1[6][24] = 4'hC;
    Number1[7][24] = 4'hC;
    Number1[8][24] = 4'hC;
    Number1[9][24] = 4'hC;
    Number1[10][24] = 4'hC;
    Number1[11][24] = 4'hC;
    Number1[12][24] = 4'hC;
    Number1[13][24] = 4'hC;
    Number1[14][24] = 4'hC;
    Number1[15][24] = 4'hC;
    Number1[16][24] = 4'hC;
    Number1[17][24] = 4'hC;
    Number1[18][24] = 4'hC;
    Number1[19][24] = 4'hC;
    Number1[20][24] = 4'hF;
    Number1[21][24] = 4'hF;
    Number1[22][24] = 4'hF;
    Number1[0][25] = 4'hF;
    Number1[1][25] = 4'hF;
    Number1[2][25] = 4'hF;
    Number1[3][25] = 4'hF;
    Number1[4][25] = 4'hD;
    Number1[5][25] = 4'hC;
    Number1[6][25] = 4'hC;
    Number1[7][25] = 4'hC;
    Number1[8][25] = 4'hC;
    Number1[9][25] = 4'hC;
    Number1[10][25] = 4'hC;
    Number1[11][25] = 4'hC;
    Number1[12][25] = 4'hC;
    Number1[13][25] = 4'hC;
    Number1[14][25] = 4'hC;
    Number1[15][25] = 4'hC;
    Number1[16][25] = 4'hC;
    Number1[17][25] = 4'hC;
    Number1[18][25] = 4'hC;
    Number1[19][25] = 4'hC;
    Number1[20][25] = 4'hF;
    Number1[21][25] = 4'hF;
    Number1[22][25] = 4'hF;
    Number1[0][26] = 4'hF;
    Number1[1][26] = 4'hF;
    Number1[2][26] = 4'hF;
    Number1[3][26] = 4'hF;
    Number1[4][26] = 4'hD;
    Number1[5][26] = 4'hC;
    Number1[6][26] = 4'hC;
    Number1[7][26] = 4'hC;
    Number1[8][26] = 4'hC;
    Number1[9][26] = 4'hC;
    Number1[10][26] = 4'hC;
    Number1[11][26] = 4'hC;
    Number1[12][26] = 4'hC;
    Number1[13][26] = 4'hC;
    Number1[14][26] = 4'hC;
    Number1[15][26] = 4'hC;
    Number1[16][26] = 4'hC;
    Number1[17][26] = 4'hC;
    Number1[18][26] = 4'hC;
    Number1[19][26] = 4'hD;
    Number1[20][26] = 4'hF;
    Number1[21][26] = 4'hF;
    Number1[22][26] = 4'hF;
    Number1[0][27] = 4'hF;
    Number1[1][27] = 4'hF;
    Number1[2][27] = 4'hF;
    Number1[3][27] = 4'hF;
    Number1[4][27] = 4'hF;
    Number1[5][27] = 4'hF;
    Number1[6][27] = 4'hF;
    Number1[7][27] = 4'hF;
    Number1[8][27] = 4'hF;
    Number1[9][27] = 4'hF;
    Number1[10][27] = 4'hF;
    Number1[11][27] = 4'hF;
    Number1[12][27] = 4'hF;
    Number1[13][27] = 4'hF;
    Number1[14][27] = 4'hF;
    Number1[15][27] = 4'hF;
    Number1[16][27] = 4'hF;
    Number1[17][27] = 4'hF;
    Number1[18][27] = 4'hF;
    Number1[19][27] = 4'hF;
    Number1[20][27] = 4'hF;
    Number1[21][27] = 4'hF;
    Number1[22][27] = 4'hF;
    Number1[0][28] = 4'hF;
    Number1[1][28] = 4'hF;
    Number1[2][28] = 4'hF;
    Number1[3][28] = 4'hF;
    Number1[4][28] = 4'hF;
    Number1[5][28] = 4'hF;
    Number1[6][28] = 4'hF;
    Number1[7][28] = 4'hF;
    Number1[8][28] = 4'hF;
    Number1[9][28] = 4'hF;
    Number1[10][28] = 4'hF;
    Number1[11][28] = 4'hF;
    Number1[12][28] = 4'hF;
    Number1[13][28] = 4'hF;
    Number1[14][28] = 4'hF;
    Number1[15][28] = 4'hF;
    Number1[16][28] = 4'hF;
    Number1[17][28] = 4'hF;
    Number1[18][28] = 4'hF;
    Number1[19][28] = 4'hF;
    Number1[20][28] = 4'hF;
    Number1[21][28] = 4'hF;
    Number1[22][28] = 4'hF;

// Number 2
    Number2[0][0] = 4'hF;
    Number2[1][0] = 4'hF;
    Number2[2][0] = 4'hF;
    Number2[3][0] = 4'hF;
    Number2[4][0] = 4'hF;
    Number2[5][0] = 4'hF;
    Number2[6][0] = 4'hF;
    Number2[7][0] = 4'hF;
    Number2[8][0] = 4'hF;
    Number2[9][0] = 4'hF;
    Number2[10][0] = 4'hF;
    Number2[11][0] = 4'hF;
    Number2[12][0] = 4'hF;
    Number2[13][0] = 4'hF;
    Number2[14][0] = 4'hF;
    Number2[15][0] = 4'hF;
    Number2[16][0] = 4'hF;
    Number2[17][0] = 4'hF;
    Number2[18][0] = 4'hF;
    Number2[19][0] = 4'hF;
    Number2[20][0] = 4'hF;
    Number2[21][0] = 4'hF;
    Number2[22][0] = 4'hF;
    Number2[0][1] = 4'hF;
    Number2[1][1] = 4'hF;
    Number2[2][1] = 4'hF;
    Number2[3][1] = 4'hF;
    Number2[4][1] = 4'hF;
    Number2[5][1] = 4'hF;
    Number2[6][1] = 4'hF;
    Number2[7][1] = 4'hF;
    Number2[8][1] = 4'hF;
    Number2[9][1] = 4'hF;
    Number2[10][1] = 4'hF;
    Number2[11][1] = 4'hF;
    Number2[12][1] = 4'hF;
    Number2[13][1] = 4'hF;
    Number2[14][1] = 4'hF;
    Number2[15][1] = 4'hF;
    Number2[16][1] = 4'hF;
    Number2[17][1] = 4'hF;
    Number2[18][1] = 4'hF;
    Number2[19][1] = 4'hF;
    Number2[20][1] = 4'hF;
    Number2[21][1] = 4'hF;
    Number2[22][1] = 4'hF;
    Number2[0][2] = 4'hF;
    Number2[1][2] = 4'hF;
    Number2[2][2] = 4'hF;
    Number2[3][2] = 4'hF;
    Number2[4][2] = 4'hF;
    Number2[5][2] = 4'hF;
    Number2[6][2] = 4'hF;
    Number2[7][2] = 4'hD;
    Number2[8][2] = 4'hD;
    Number2[9][2] = 4'hC;
    Number2[10][2] = 4'hC;
    Number2[11][2] = 4'hC;
    Number2[12][2] = 4'hC;
    Number2[13][2] = 4'hC;
    Number2[14][2] = 4'hD;
    Number2[15][2] = 4'hE;
    Number2[16][2] = 4'hF;
    Number2[17][2] = 4'hF;
    Number2[18][2] = 4'hF;
    Number2[19][2] = 4'hF;
    Number2[20][2] = 4'hF;
    Number2[21][2] = 4'hF;
    Number2[22][2] = 4'hF;
    Number2[0][3] = 4'hF;
    Number2[1][3] = 4'hF;
    Number2[2][3] = 4'hF;
    Number2[3][3] = 4'hF;
    Number2[4][3] = 4'hF;
    Number2[5][3] = 4'hD;
    Number2[6][3] = 4'hC;
    Number2[7][3] = 4'hC;
    Number2[8][3] = 4'hC;
    Number2[9][3] = 4'hC;
    Number2[10][3] = 4'hC;
    Number2[11][3] = 4'hC;
    Number2[12][3] = 4'hC;
    Number2[13][3] = 4'hC;
    Number2[14][3] = 4'hC;
    Number2[15][3] = 4'hC;
    Number2[16][3] = 4'hD;
    Number2[17][3] = 4'hE;
    Number2[18][3] = 4'hF;
    Number2[19][3] = 4'hF;
    Number2[20][3] = 4'hF;
    Number2[21][3] = 4'hF;
    Number2[22][3] = 4'hF;
    Number2[0][4] = 4'hF;
    Number2[1][4] = 4'hF;
    Number2[2][4] = 4'hF;
    Number2[3][4] = 4'hE;
    Number2[4][4] = 4'hC;
    Number2[5][4] = 4'hC;
    Number2[6][4] = 4'hC;
    Number2[7][4] = 4'hC;
    Number2[8][4] = 4'hC;
    Number2[9][4] = 4'hC;
    Number2[10][4] = 4'hC;
    Number2[11][4] = 4'hC;
    Number2[12][4] = 4'hC;
    Number2[13][4] = 4'hC;
    Number2[14][4] = 4'hC;
    Number2[15][4] = 4'hC;
    Number2[16][4] = 4'hC;
    Number2[17][4] = 4'hC;
    Number2[18][4] = 4'hF;
    Number2[19][4] = 4'hF;
    Number2[20][4] = 4'hF;
    Number2[21][4] = 4'hF;
    Number2[22][4] = 4'hF;
    Number2[0][5] = 4'hF;
    Number2[1][5] = 4'hF;
    Number2[2][5] = 4'hF;
    Number2[3][5] = 4'hD;
    Number2[4][5] = 4'hC;
    Number2[5][5] = 4'hC;
    Number2[6][5] = 4'hC;
    Number2[7][5] = 4'hC;
    Number2[8][5] = 4'hC;
    Number2[9][5] = 4'hC;
    Number2[10][5] = 4'hC;
    Number2[11][5] = 4'hC;
    Number2[12][5] = 4'hC;
    Number2[13][5] = 4'hC;
    Number2[14][5] = 4'hC;
    Number2[15][5] = 4'hC;
    Number2[16][5] = 4'hC;
    Number2[17][5] = 4'hC;
    Number2[18][5] = 4'hD;
    Number2[19][5] = 4'hF;
    Number2[20][5] = 4'hF;
    Number2[21][5] = 4'hF;
    Number2[22][5] = 4'hF;
    Number2[0][6] = 4'hF;
    Number2[1][6] = 4'hF;
    Number2[2][6] = 4'hF;
    Number2[3][6] = 4'hD;
    Number2[4][6] = 4'hC;
    Number2[5][6] = 4'hC;
    Number2[6][6] = 4'hC;
    Number2[7][6] = 4'hD;
    Number2[8][6] = 4'hE;
    Number2[9][6] = 4'hF;
    Number2[10][6] = 4'hE;
    Number2[11][6] = 4'hD;
    Number2[12][6] = 4'hC;
    Number2[13][6] = 4'hC;
    Number2[14][6] = 4'hC;
    Number2[15][6] = 4'hC;
    Number2[16][6] = 4'hC;
    Number2[17][6] = 4'hC;
    Number2[18][6] = 4'hC;
    Number2[19][6] = 4'hF;
    Number2[20][6] = 4'hF;
    Number2[21][6] = 4'hF;
    Number2[22][6] = 4'hF;
    Number2[0][7] = 4'hF;
    Number2[1][7] = 4'hF;
    Number2[2][7] = 4'hF;
    Number2[3][7] = 4'hE;
    Number2[4][7] = 4'hC;
    Number2[5][7] = 4'hD;
    Number2[6][7] = 4'hF;
    Number2[7][7] = 4'hF;
    Number2[8][7] = 4'hF;
    Number2[9][7] = 4'hF;
    Number2[10][7] = 4'hF;
    Number2[11][7] = 4'hF;
    Number2[12][7] = 4'hD;
    Number2[13][7] = 4'hC;
    Number2[14][7] = 4'hC;
    Number2[15][7] = 4'hC;
    Number2[16][7] = 4'hC;
    Number2[17][7] = 4'hC;
    Number2[18][7] = 4'hC;
    Number2[19][7] = 4'hE;
    Number2[20][7] = 4'hF;
    Number2[21][7] = 4'hF;
    Number2[22][7] = 4'hF;
    Number2[0][8] = 4'hF;
    Number2[1][8] = 4'hF;
    Number2[2][8] = 4'hF;
    Number2[3][8] = 4'hF;
    Number2[4][8] = 4'hF;
    Number2[5][8] = 4'hF;
    Number2[6][8] = 4'hF;
    Number2[7][8] = 4'hF;
    Number2[8][8] = 4'hF;
    Number2[9][8] = 4'hF;
    Number2[10][8] = 4'hF;
    Number2[11][8] = 4'hF;
    Number2[12][8] = 4'hE;
    Number2[13][8] = 4'hC;
    Number2[14][8] = 4'hC;
    Number2[15][8] = 4'hC;
    Number2[16][8] = 4'hC;
    Number2[17][8] = 4'hC;
    Number2[18][8] = 4'hC;
    Number2[19][8] = 4'hE;
    Number2[20][8] = 4'hF;
    Number2[21][8] = 4'hF;
    Number2[22][8] = 4'hF;
    Number2[0][9] = 4'hF;
    Number2[1][9] = 4'hF;
    Number2[2][9] = 4'hF;
    Number2[3][9] = 4'hF;
    Number2[4][9] = 4'hF;
    Number2[5][9] = 4'hF;
    Number2[6][9] = 4'hF;
    Number2[7][9] = 4'hF;
    Number2[8][9] = 4'hF;
    Number2[9][9] = 4'hF;
    Number2[10][9] = 4'hF;
    Number2[11][9] = 4'hF;
    Number2[12][9] = 4'hF;
    Number2[13][9] = 4'hC;
    Number2[14][9] = 4'hC;
    Number2[15][9] = 4'hC;
    Number2[16][9] = 4'hC;
    Number2[17][9] = 4'hC;
    Number2[18][9] = 4'hC;
    Number2[19][9] = 4'hF;
    Number2[20][9] = 4'hF;
    Number2[21][9] = 4'hF;
    Number2[22][9] = 4'hF;
    Number2[0][10] = 4'hF;
    Number2[1][10] = 4'hF;
    Number2[2][10] = 4'hF;
    Number2[3][10] = 4'hF;
    Number2[4][10] = 4'hF;
    Number2[5][10] = 4'hF;
    Number2[6][10] = 4'hF;
    Number2[7][10] = 4'hF;
    Number2[8][10] = 4'hF;
    Number2[9][10] = 4'hF;
    Number2[10][10] = 4'hF;
    Number2[11][10] = 4'hF;
    Number2[12][10] = 4'hE;
    Number2[13][10] = 4'hC;
    Number2[14][10] = 4'hC;
    Number2[15][10] = 4'hC;
    Number2[16][10] = 4'hC;
    Number2[17][10] = 4'hC;
    Number2[18][10] = 4'hC;
    Number2[19][10] = 4'hF;
    Number2[20][10] = 4'hF;
    Number2[21][10] = 4'hF;
    Number2[22][10] = 4'hF;
    Number2[0][11] = 4'hF;
    Number2[1][11] = 4'hF;
    Number2[2][11] = 4'hF;
    Number2[3][11] = 4'hF;
    Number2[4][11] = 4'hF;
    Number2[5][11] = 4'hF;
    Number2[6][11] = 4'hF;
    Number2[7][11] = 4'hF;
    Number2[8][11] = 4'hF;
    Number2[9][11] = 4'hF;
    Number2[10][11] = 4'hF;
    Number2[11][11] = 4'hF;
    Number2[12][11] = 4'hD;
    Number2[13][11] = 4'hC;
    Number2[14][11] = 4'hC;
    Number2[15][11] = 4'hC;
    Number2[16][11] = 4'hC;
    Number2[17][11] = 4'hC;
    Number2[18][11] = 4'hC;
    Number2[19][11] = 4'hF;
    Number2[20][11] = 4'hF;
    Number2[21][11] = 4'hF;
    Number2[22][11] = 4'hF;
    Number2[0][12] = 4'hF;
    Number2[1][12] = 4'hF;
    Number2[2][12] = 4'hF;
    Number2[3][12] = 4'hF;
    Number2[4][12] = 4'hF;
    Number2[5][12] = 4'hF;
    Number2[6][12] = 4'hF;
    Number2[7][12] = 4'hF;
    Number2[8][12] = 4'hF;
    Number2[9][12] = 4'hF;
    Number2[10][12] = 4'hF;
    Number2[11][12] = 4'hF;
    Number2[12][12] = 4'hD;
    Number2[13][12] = 4'hC;
    Number2[14][12] = 4'hC;
    Number2[15][12] = 4'hC;
    Number2[16][12] = 4'hC;
    Number2[17][12] = 4'hC;
    Number2[18][12] = 4'hD;
    Number2[19][12] = 4'hF;
    Number2[20][12] = 4'hF;
    Number2[21][12] = 4'hF;
    Number2[22][12] = 4'hF;
    Number2[0][13] = 4'hF;
    Number2[1][13] = 4'hF;
    Number2[2][13] = 4'hF;
    Number2[3][13] = 4'hF;
    Number2[4][13] = 4'hF;
    Number2[5][13] = 4'hF;
    Number2[6][13] = 4'hF;
    Number2[7][13] = 4'hF;
    Number2[8][13] = 4'hF;
    Number2[9][13] = 4'hF;
    Number2[10][13] = 4'hF;
    Number2[11][13] = 4'hD;
    Number2[12][13] = 4'hC;
    Number2[13][13] = 4'hC;
    Number2[14][13] = 4'hC;
    Number2[15][13] = 4'hC;
    Number2[16][13] = 4'hC;
    Number2[17][13] = 4'hC;
    Number2[18][13] = 4'hF;
    Number2[19][13] = 4'hF;
    Number2[20][13] = 4'hF;
    Number2[21][13] = 4'hF;
    Number2[22][13] = 4'hF;
    Number2[0][14] = 4'hF;
    Number2[1][14] = 4'hF;
    Number2[2][14] = 4'hF;
    Number2[3][14] = 4'hF;
    Number2[4][14] = 4'hF;
    Number2[5][14] = 4'hF;
    Number2[6][14] = 4'hF;
    Number2[7][14] = 4'hF;
    Number2[8][14] = 4'hF;
    Number2[9][14] = 4'hF;
    Number2[10][14] = 4'hE;
    Number2[11][14] = 4'hC;
    Number2[12][14] = 4'hC;
    Number2[13][14] = 4'hC;
    Number2[14][14] = 4'hC;
    Number2[15][14] = 4'hC;
    Number2[16][14] = 4'hC;
    Number2[17][14] = 4'hE;
    Number2[18][14] = 4'hF;
    Number2[19][14] = 4'hF;
    Number2[20][14] = 4'hF;
    Number2[21][14] = 4'hF;
    Number2[22][14] = 4'hF;
    Number2[0][15] = 4'hF;
    Number2[1][15] = 4'hF;
    Number2[2][15] = 4'hF;
    Number2[3][15] = 4'hF;
    Number2[4][15] = 4'hF;
    Number2[5][15] = 4'hF;
    Number2[6][15] = 4'hF;
    Number2[7][15] = 4'hF;
    Number2[8][15] = 4'hF;
    Number2[9][15] = 4'hF;
    Number2[10][15] = 4'hC;
    Number2[11][15] = 4'hC;
    Number2[12][15] = 4'hC;
    Number2[13][15] = 4'hC;
    Number2[14][15] = 4'hC;
    Number2[15][15] = 4'hC;
    Number2[16][15] = 4'hD;
    Number2[17][15] = 4'hF;
    Number2[18][15] = 4'hF;
    Number2[19][15] = 4'hF;
    Number2[20][15] = 4'hF;
    Number2[21][15] = 4'hF;
    Number2[22][15] = 4'hF;
    Number2[0][16] = 4'hF;
    Number2[1][16] = 4'hF;
    Number2[2][16] = 4'hF;
    Number2[3][16] = 4'hF;
    Number2[4][16] = 4'hF;
    Number2[5][16] = 4'hF;
    Number2[6][16] = 4'hF;
    Number2[7][16] = 4'hF;
    Number2[8][16] = 4'hF;
    Number2[9][16] = 4'hD;
    Number2[10][16] = 4'hC;
    Number2[11][16] = 4'hC;
    Number2[12][16] = 4'hC;
    Number2[13][16] = 4'hC;
    Number2[14][16] = 4'hC;
    Number2[15][16] = 4'hD;
    Number2[16][16] = 4'hF;
    Number2[17][16] = 4'hF;
    Number2[18][16] = 4'hF;
    Number2[19][16] = 4'hF;
    Number2[20][16] = 4'hF;
    Number2[21][16] = 4'hF;
    Number2[22][16] = 4'hF;
    Number2[0][17] = 4'hF;
    Number2[1][17] = 4'hF;
    Number2[2][17] = 4'hF;
    Number2[3][17] = 4'hF;
    Number2[4][17] = 4'hF;
    Number2[5][17] = 4'hF;
    Number2[6][17] = 4'hF;
    Number2[7][17] = 4'hF;
    Number2[8][17] = 4'hD;
    Number2[9][17] = 4'hC;
    Number2[10][17] = 4'hC;
    Number2[11][17] = 4'hC;
    Number2[12][17] = 4'hC;
    Number2[13][17] = 4'hC;
    Number2[14][17] = 4'hD;
    Number2[15][17] = 4'hF;
    Number2[16][17] = 4'hF;
    Number2[17][17] = 4'hF;
    Number2[18][17] = 4'hF;
    Number2[19][17] = 4'hF;
    Number2[20][17] = 4'hF;
    Number2[21][17] = 4'hF;
    Number2[22][17] = 4'hF;
    Number2[0][18] = 4'hF;
    Number2[1][18] = 4'hF;
    Number2[2][18] = 4'hF;
    Number2[3][18] = 4'hF;
    Number2[4][18] = 4'hF;
    Number2[5][18] = 4'hF;
    Number2[6][18] = 4'hF;
    Number2[7][18] = 4'hD;
    Number2[8][18] = 4'hC;
    Number2[9][18] = 4'hC;
    Number2[10][18] = 4'hC;
    Number2[11][18] = 4'hC;
    Number2[12][18] = 4'hC;
    Number2[13][18] = 4'hC;
    Number2[14][18] = 4'hF;
    Number2[15][18] = 4'hF;
    Number2[16][18] = 4'hF;
    Number2[17][18] = 4'hF;
    Number2[18][18] = 4'hF;
    Number2[19][18] = 4'hF;
    Number2[20][18] = 4'hF;
    Number2[21][18] = 4'hF;
    Number2[22][18] = 4'hF;
    Number2[0][19] = 4'hF;
    Number2[1][19] = 4'hF;
    Number2[2][19] = 4'hF;
    Number2[3][19] = 4'hF;
    Number2[4][19] = 4'hF;
    Number2[5][19] = 4'hF;
    Number2[6][19] = 4'hD;
    Number2[7][19] = 4'hC;
    Number2[8][19] = 4'hC;
    Number2[9][19] = 4'hC;
    Number2[10][19] = 4'hC;
    Number2[11][19] = 4'hC;
    Number2[12][19] = 4'hC;
    Number2[13][19] = 4'hF;
    Number2[14][19] = 4'hF;
    Number2[15][19] = 4'hF;
    Number2[16][19] = 4'hF;
    Number2[17][19] = 4'hF;
    Number2[18][19] = 4'hF;
    Number2[19][19] = 4'hF;
    Number2[20][19] = 4'hF;
    Number2[21][19] = 4'hF;
    Number2[22][19] = 4'hF;
    Number2[0][20] = 4'hF;
    Number2[1][20] = 4'hF;
    Number2[2][20] = 4'hF;
    Number2[3][20] = 4'hF;
    Number2[4][20] = 4'hF;
    Number2[5][20] = 4'hD;
    Number2[6][20] = 4'hC;
    Number2[7][20] = 4'hC;
    Number2[8][20] = 4'hC;
    Number2[9][20] = 4'hC;
    Number2[10][20] = 4'hC;
    Number2[11][20] = 4'hC;
    Number2[12][20] = 4'hF;
    Number2[13][20] = 4'hF;
    Number2[14][20] = 4'hF;
    Number2[15][20] = 4'hF;
    Number2[16][20] = 4'hF;
    Number2[17][20] = 4'hF;
    Number2[18][20] = 4'hF;
    Number2[19][20] = 4'hF;
    Number2[20][20] = 4'hF;
    Number2[21][20] = 4'hF;
    Number2[22][20] = 4'hF;
    Number2[0][21] = 4'hF;
    Number2[1][21] = 4'hF;
    Number2[2][21] = 4'hF;
    Number2[3][21] = 4'hF;
    Number2[4][21] = 4'hD;
    Number2[5][21] = 4'hC;
    Number2[6][21] = 4'hC;
    Number2[7][21] = 4'hC;
    Number2[8][21] = 4'hC;
    Number2[9][21] = 4'hC;
    Number2[10][21] = 4'hC;
    Number2[11][21] = 4'hF;
    Number2[12][21] = 4'hF;
    Number2[13][21] = 4'hF;
    Number2[14][21] = 4'hF;
    Number2[15][21] = 4'hF;
    Number2[16][21] = 4'hF;
    Number2[17][21] = 4'hF;
    Number2[18][21] = 4'hF;
    Number2[19][21] = 4'hF;
    Number2[20][21] = 4'hF;
    Number2[21][21] = 4'hF;
    Number2[22][21] = 4'hF;
    Number2[0][22] = 4'hF;
    Number2[1][22] = 4'hF;
    Number2[2][22] = 4'hF;
    Number2[3][22] = 4'hE;
    Number2[4][22] = 4'hC;
    Number2[5][22] = 4'hC;
    Number2[6][22] = 4'hC;
    Number2[7][22] = 4'hC;
    Number2[8][22] = 4'hC;
    Number2[9][22] = 4'hC;
    Number2[10][22] = 4'hF;
    Number2[11][22] = 4'hF;
    Number2[12][22] = 4'hF;
    Number2[13][22] = 4'hF;
    Number2[14][22] = 4'hF;
    Number2[15][22] = 4'hF;
    Number2[16][22] = 4'hF;
    Number2[17][22] = 4'hF;
    Number2[18][22] = 4'hF;
    Number2[19][22] = 4'hF;
    Number2[20][22] = 4'hF;
    Number2[21][22] = 4'hF;
    Number2[22][22] = 4'hF;
    Number2[0][23] = 4'hF;
    Number2[1][23] = 4'hF;
    Number2[2][23] = 4'hF;
    Number2[3][23] = 4'hD;
    Number2[4][23] = 4'hC;
    Number2[5][23] = 4'hC;
    Number2[6][23] = 4'hC;
    Number2[7][23] = 4'hC;
    Number2[8][23] = 4'hC;
    Number2[9][23] = 4'hC;
    Number2[10][23] = 4'hC;
    Number2[11][23] = 4'hC;
    Number2[12][23] = 4'hC;
    Number2[13][23] = 4'hC;
    Number2[14][23] = 4'hC;
    Number2[15][23] = 4'hC;
    Number2[16][23] = 4'hC;
    Number2[17][23] = 4'hC;
    Number2[18][23] = 4'hC;
    Number2[19][23] = 4'hC;
    Number2[20][23] = 4'hF;
    Number2[21][23] = 4'hF;
    Number2[22][23] = 4'hF;
    Number2[0][24] = 4'hF;
    Number2[1][24] = 4'hF;
    Number2[2][24] = 4'hF;
    Number2[3][24] = 4'hC;
    Number2[4][24] = 4'hC;
    Number2[5][24] = 4'hC;
    Number2[6][24] = 4'hC;
    Number2[7][24] = 4'hC;
    Number2[8][24] = 4'hC;
    Number2[9][24] = 4'hC;
    Number2[10][24] = 4'hC;
    Number2[11][24] = 4'hC;
    Number2[12][24] = 4'hC;
    Number2[13][24] = 4'hC;
    Number2[14][24] = 4'hC;
    Number2[15][24] = 4'hC;
    Number2[16][24] = 4'hC;
    Number2[17][24] = 4'hC;
    Number2[18][24] = 4'hC;
    Number2[19][24] = 4'hC;
    Number2[20][24] = 4'hE;
    Number2[21][24] = 4'hF;
    Number2[22][24] = 4'hF;
    Number2[0][25] = 4'hF;
    Number2[1][25] = 4'hF;
    Number2[2][25] = 4'hF;
    Number2[3][25] = 4'hC;
    Number2[4][25] = 4'hC;
    Number2[5][25] = 4'hC;
    Number2[6][25] = 4'hC;
    Number2[7][25] = 4'hC;
    Number2[8][25] = 4'hC;
    Number2[9][25] = 4'hC;
    Number2[10][25] = 4'hC;
    Number2[11][25] = 4'hC;
    Number2[12][25] = 4'hC;
    Number2[13][25] = 4'hC;
    Number2[14][25] = 4'hC;
    Number2[15][25] = 4'hC;
    Number2[16][25] = 4'hC;
    Number2[17][25] = 4'hC;
    Number2[18][25] = 4'hC;
    Number2[19][25] = 4'hC;
    Number2[20][25] = 4'hE;
    Number2[21][25] = 4'hF;
    Number2[22][25] = 4'hF;
    Number2[0][26] = 4'hF;
    Number2[1][26] = 4'hF;
    Number2[2][26] = 4'hF;
    Number2[3][26] = 4'hD;
    Number2[4][26] = 4'hC;
    Number2[5][26] = 4'hC;
    Number2[6][26] = 4'hC;
    Number2[7][26] = 4'hC;
    Number2[8][26] = 4'hC;
    Number2[9][26] = 4'hC;
    Number2[10][26] = 4'hC;
    Number2[11][26] = 4'hC;
    Number2[12][26] = 4'hC;
    Number2[13][26] = 4'hC;
    Number2[14][26] = 4'hC;
    Number2[15][26] = 4'hC;
    Number2[16][26] = 4'hC;
    Number2[17][26] = 4'hC;
    Number2[18][26] = 4'hC;
    Number2[19][26] = 4'hC;
    Number2[20][26] = 4'hF;
    Number2[21][26] = 4'hF;
    Number2[22][26] = 4'hF;
    Number2[0][27] = 4'hF;
    Number2[1][27] = 4'hF;
    Number2[2][27] = 4'hF;
    Number2[3][27] = 4'hF;
    Number2[4][27] = 4'hF;
    Number2[5][27] = 4'hF;
    Number2[6][27] = 4'hF;
    Number2[7][27] = 4'hF;
    Number2[8][27] = 4'hF;
    Number2[9][27] = 4'hF;
    Number2[10][27] = 4'hF;
    Number2[11][27] = 4'hF;
    Number2[12][27] = 4'hF;
    Number2[13][27] = 4'hF;
    Number2[14][27] = 4'hF;
    Number2[15][27] = 4'hF;
    Number2[16][27] = 4'hF;
    Number2[17][27] = 4'hF;
    Number2[18][27] = 4'hF;
    Number2[19][27] = 4'hF;
    Number2[20][27] = 4'hF;
    Number2[21][27] = 4'hF;
    Number2[22][27] = 4'hF;
    Number2[0][28] = 4'hF;
    Number2[1][28] = 4'hF;
    Number2[2][28] = 4'hF;
    Number2[3][28] = 4'hF;
    Number2[4][28] = 4'hF;
    Number2[5][28] = 4'hF;
    Number2[6][28] = 4'hF;
    Number2[7][28] = 4'hF;
    Number2[8][28] = 4'hF;
    Number2[9][28] = 4'hF;
    Number2[10][28] = 4'hF;
    Number2[11][28] = 4'hF;
    Number2[12][28] = 4'hF;
    Number2[13][28] = 4'hF;
    Number2[14][28] = 4'hF;
    Number2[15][28] = 4'hF;
    Number2[16][28] = 4'hF;
    Number2[17][28] = 4'hF;
    Number2[18][28] = 4'hF;
    Number2[19][28] = 4'hF;
    Number2[20][28] = 4'hF;
    Number2[21][28] = 4'hF;
    Number2[22][28] = 4'hF;

// Number 3
    Number3[0][0] = 4'hF;
    Number3[1][0] = 4'hF;
    Number3[2][0] = 4'hF;
    Number3[3][0] = 4'hF;
    Number3[4][0] = 4'hF;
    Number3[5][0] = 4'hF;
    Number3[6][0] = 4'hF;
    Number3[7][0] = 4'hF;
    Number3[8][0] = 4'hF;
    Number3[9][0] = 4'hF;
    Number3[10][0] = 4'hF;
    Number3[11][0] = 4'hF;
    Number3[12][0] = 4'hF;
    Number3[13][0] = 4'hF;
    Number3[14][0] = 4'hF;
    Number3[15][0] = 4'hF;
    Number3[16][0] = 4'hF;
    Number3[17][0] = 4'hF;
    Number3[18][0] = 4'hF;
    Number3[19][0] = 4'hF;
    Number3[20][0] = 4'hF;
    Number3[21][0] = 4'hF;
    Number3[22][0] = 4'hF;
    Number3[0][1] = 4'hF;
    Number3[1][1] = 4'hF;
    Number3[2][1] = 4'hF;
    Number3[3][1] = 4'hF;
    Number3[4][1] = 4'hF;
    Number3[5][1] = 4'hF;
    Number3[6][1] = 4'hF;
    Number3[7][1] = 4'hF;
    Number3[8][1] = 4'hF;
    Number3[9][1] = 4'hF;
    Number3[10][1] = 4'hF;
    Number3[11][1] = 4'hF;
    Number3[12][1] = 4'hF;
    Number3[13][1] = 4'hF;
    Number3[14][1] = 4'hF;
    Number3[15][1] = 4'hF;
    Number3[16][1] = 4'hF;
    Number3[17][1] = 4'hF;
    Number3[18][1] = 4'hF;
    Number3[19][1] = 4'hF;
    Number3[20][1] = 4'hF;
    Number3[21][1] = 4'hF;
    Number3[22][1] = 4'hF;
    Number3[0][2] = 4'hF;
    Number3[1][2] = 4'hF;
    Number3[2][2] = 4'hF;
    Number3[3][2] = 4'hF;
    Number3[4][2] = 4'hF;
    Number3[5][2] = 4'hF;
    Number3[6][2] = 4'hE;
    Number3[7][2] = 4'hD;
    Number3[8][2] = 4'hD;
    Number3[9][2] = 4'hC;
    Number3[10][2] = 4'hC;
    Number3[11][2] = 4'hC;
    Number3[12][2] = 4'hC;
    Number3[13][2] = 4'hC;
    Number3[14][2] = 4'hD;
    Number3[15][2] = 4'hE;
    Number3[16][2] = 4'hF;
    Number3[17][2] = 4'hF;
    Number3[18][2] = 4'hF;
    Number3[19][2] = 4'hF;
    Number3[20][2] = 4'hF;
    Number3[21][2] = 4'hF;
    Number3[22][2] = 4'hF;
    Number3[0][3] = 4'hF;
    Number3[1][3] = 4'hF;
    Number3[2][3] = 4'hF;
    Number3[3][3] = 4'hF;
    Number3[4][3] = 4'hE;
    Number3[5][3] = 4'hD;
    Number3[6][3] = 4'hC;
    Number3[7][3] = 4'hC;
    Number3[8][3] = 4'hC;
    Number3[9][3] = 4'hC;
    Number3[10][3] = 4'hC;
    Number3[11][3] = 4'hC;
    Number3[12][3] = 4'hC;
    Number3[13][3] = 4'hC;
    Number3[14][3] = 4'hC;
    Number3[15][3] = 4'hC;
    Number3[16][3] = 4'hC;
    Number3[17][3] = 4'hE;
    Number3[18][3] = 4'hF;
    Number3[19][3] = 4'hF;
    Number3[20][3] = 4'hF;
    Number3[21][3] = 4'hF;
    Number3[22][3] = 4'hF;
    Number3[0][4] = 4'hF;
    Number3[1][4] = 4'hF;
    Number3[2][4] = 4'hF;
    Number3[3][4] = 4'hE;
    Number3[4][4] = 4'hC;
    Number3[5][4] = 4'hC;
    Number3[6][4] = 4'hC;
    Number3[7][4] = 4'hC;
    Number3[8][4] = 4'hC;
    Number3[9][4] = 4'hC;
    Number3[10][4] = 4'hC;
    Number3[11][4] = 4'hC;
    Number3[12][4] = 4'hC;
    Number3[13][4] = 4'hC;
    Number3[14][4] = 4'hC;
    Number3[15][4] = 4'hC;
    Number3[16][4] = 4'hC;
    Number3[17][4] = 4'hC;
    Number3[18][4] = 4'hF;
    Number3[19][4] = 4'hF;
    Number3[20][4] = 4'hF;
    Number3[21][4] = 4'hF;
    Number3[22][4] = 4'hF;
    Number3[0][5] = 4'hF;
    Number3[1][5] = 4'hF;
    Number3[2][5] = 4'hF;
    Number3[3][5] = 4'hE;
    Number3[4][5] = 4'hC;
    Number3[5][5] = 4'hC;
    Number3[6][5] = 4'hC;
    Number3[7][5] = 4'hC;
    Number3[8][5] = 4'hC;
    Number3[9][5] = 4'hC;
    Number3[10][5] = 4'hC;
    Number3[11][5] = 4'hC;
    Number3[12][5] = 4'hC;
    Number3[13][5] = 4'hC;
    Number3[14][5] = 4'hC;
    Number3[15][5] = 4'hC;
    Number3[16][5] = 4'hC;
    Number3[17][5] = 4'hC;
    Number3[18][5] = 4'hD;
    Number3[19][5] = 4'hF;
    Number3[20][5] = 4'hF;
    Number3[21][5] = 4'hF;
    Number3[22][5] = 4'hF;
    Number3[0][6] = 4'hF;
    Number3[1][6] = 4'hF;
    Number3[2][6] = 4'hF;
    Number3[3][6] = 4'hD;
    Number3[4][6] = 4'hC;
    Number3[5][6] = 4'hC;
    Number3[6][6] = 4'hC;
    Number3[7][6] = 4'hD;
    Number3[8][6] = 4'hE;
    Number3[9][6] = 4'hF;
    Number3[10][6] = 4'hE;
    Number3[11][6] = 4'hD;
    Number3[12][6] = 4'hC;
    Number3[13][6] = 4'hC;
    Number3[14][6] = 4'hC;
    Number3[15][6] = 4'hC;
    Number3[16][6] = 4'hC;
    Number3[17][6] = 4'hC;
    Number3[18][6] = 4'hC;
    Number3[19][6] = 4'hF;
    Number3[20][6] = 4'hF;
    Number3[21][6] = 4'hF;
    Number3[22][6] = 4'hF;
    Number3[0][7] = 4'hF;
    Number3[1][7] = 4'hF;
    Number3[2][7] = 4'hF;
    Number3[3][7] = 4'hE;
    Number3[4][7] = 4'hC;
    Number3[5][7] = 4'hD;
    Number3[6][7] = 4'hF;
    Number3[7][7] = 4'hF;
    Number3[8][7] = 4'hF;
    Number3[9][7] = 4'hF;
    Number3[10][7] = 4'hF;
    Number3[11][7] = 4'hF;
    Number3[12][7] = 4'hE;
    Number3[13][7] = 4'hC;
    Number3[14][7] = 4'hC;
    Number3[15][7] = 4'hC;
    Number3[16][7] = 4'hC;
    Number3[17][7] = 4'hC;
    Number3[18][7] = 4'hC;
    Number3[19][7] = 4'hF;
    Number3[20][7] = 4'hF;
    Number3[21][7] = 4'hF;
    Number3[22][7] = 4'hF;
    Number3[0][8] = 4'hF;
    Number3[1][8] = 4'hF;
    Number3[2][8] = 4'hF;
    Number3[3][8] = 4'hF;
    Number3[4][8] = 4'hF;
    Number3[5][8] = 4'hF;
    Number3[6][8] = 4'hF;
    Number3[7][8] = 4'hF;
    Number3[8][8] = 4'hF;
    Number3[9][8] = 4'hF;
    Number3[10][8] = 4'hF;
    Number3[11][8] = 4'hF;
    Number3[12][8] = 4'hF;
    Number3[13][8] = 4'hC;
    Number3[14][8] = 4'hC;
    Number3[15][8] = 4'hC;
    Number3[16][8] = 4'hC;
    Number3[17][8] = 4'hC;
    Number3[18][8] = 4'hC;
    Number3[19][8] = 4'hF;
    Number3[20][8] = 4'hF;
    Number3[21][8] = 4'hF;
    Number3[22][8] = 4'hF;
    Number3[0][9] = 4'hF;
    Number3[1][9] = 4'hF;
    Number3[2][9] = 4'hF;
    Number3[3][9] = 4'hF;
    Number3[4][9] = 4'hF;
    Number3[5][9] = 4'hF;
    Number3[6][9] = 4'hF;
    Number3[7][9] = 4'hF;
    Number3[8][9] = 4'hF;
    Number3[9][9] = 4'hF;
    Number3[10][9] = 4'hF;
    Number3[11][9] = 4'hF;
    Number3[12][9] = 4'hF;
    Number3[13][9] = 4'hC;
    Number3[14][9] = 4'hC;
    Number3[15][9] = 4'hC;
    Number3[16][9] = 4'hC;
    Number3[17][9] = 4'hC;
    Number3[18][9] = 4'hC;
    Number3[19][9] = 4'hF;
    Number3[20][9] = 4'hF;
    Number3[21][9] = 4'hF;
    Number3[22][9] = 4'hF;
    Number3[0][10] = 4'hF;
    Number3[1][10] = 4'hF;
    Number3[2][10] = 4'hF;
    Number3[3][10] = 4'hF;
    Number3[4][10] = 4'hF;
    Number3[5][10] = 4'hF;
    Number3[6][10] = 4'hF;
    Number3[7][10] = 4'hF;
    Number3[8][10] = 4'hF;
    Number3[9][10] = 4'hF;
    Number3[10][10] = 4'hF;
    Number3[11][10] = 4'hF;
    Number3[12][10] = 4'hD;
    Number3[13][10] = 4'hC;
    Number3[14][10] = 4'hC;
    Number3[15][10] = 4'hC;
    Number3[16][10] = 4'hC;
    Number3[17][10] = 4'hC;
    Number3[18][10] = 4'hD;
    Number3[19][10] = 4'hF;
    Number3[20][10] = 4'hF;
    Number3[21][10] = 4'hF;
    Number3[22][10] = 4'hF;
    Number3[0][11] = 4'hF;
    Number3[1][11] = 4'hF;
    Number3[2][11] = 4'hF;
    Number3[3][11] = 4'hF;
    Number3[4][11] = 4'hF;
    Number3[5][11] = 4'hF;
    Number3[6][11] = 4'hF;
    Number3[7][11] = 4'hF;
    Number3[8][11] = 4'hF;
    Number3[9][11] = 4'hF;
    Number3[10][11] = 4'hE;
    Number3[11][11] = 4'hD;
    Number3[12][11] = 4'hC;
    Number3[13][11] = 4'hC;
    Number3[14][11] = 4'hC;
    Number3[15][11] = 4'hC;
    Number3[16][11] = 4'hC;
    Number3[17][11] = 4'hC;
    Number3[18][11] = 4'hF;
    Number3[19][11] = 4'hF;
    Number3[20][11] = 4'hF;
    Number3[21][11] = 4'hF;
    Number3[22][11] = 4'hF;
    Number3[0][12] = 4'hF;
    Number3[1][12] = 4'hF;
    Number3[2][12] = 4'hF;
    Number3[3][12] = 4'hF;
    Number3[4][12] = 4'hF;
    Number3[5][12] = 4'hD;
    Number3[6][12] = 4'hC;
    Number3[7][12] = 4'hC;
    Number3[8][12] = 4'hC;
    Number3[9][12] = 4'hC;
    Number3[10][12] = 4'hC;
    Number3[11][12] = 4'hC;
    Number3[12][12] = 4'hC;
    Number3[13][12] = 4'hC;
    Number3[14][12] = 4'hC;
    Number3[15][12] = 4'hC;
    Number3[16][12] = 4'hD;
    Number3[17][12] = 4'hF;
    Number3[18][12] = 4'hF;
    Number3[19][12] = 4'hF;
    Number3[20][12] = 4'hF;
    Number3[21][12] = 4'hF;
    Number3[22][12] = 4'hF;
    Number3[0][13] = 4'hF;
    Number3[1][13] = 4'hF;
    Number3[2][13] = 4'hF;
    Number3[3][13] = 4'hF;
    Number3[4][13] = 4'hF;
    Number3[5][13] = 4'hD;
    Number3[6][13] = 4'hC;
    Number3[7][13] = 4'hC;
    Number3[8][13] = 4'hC;
    Number3[9][13] = 4'hC;
    Number3[10][13] = 4'hC;
    Number3[11][13] = 4'hC;
    Number3[12][13] = 4'hC;
    Number3[13][13] = 4'hC;
    Number3[14][13] = 4'hC;
    Number3[15][13] = 4'hD;
    Number3[16][13] = 4'hF;
    Number3[17][13] = 4'hF;
    Number3[18][13] = 4'hF;
    Number3[19][13] = 4'hF;
    Number3[20][13] = 4'hF;
    Number3[21][13] = 4'hF;
    Number3[22][13] = 4'hF;
    Number3[0][14] = 4'hF;
    Number3[1][14] = 4'hF;
    Number3[2][14] = 4'hF;
    Number3[3][14] = 4'hF;
    Number3[4][14] = 4'hF;
    Number3[5][14] = 4'hD;
    Number3[6][14] = 4'hC;
    Number3[7][14] = 4'hC;
    Number3[8][14] = 4'hC;
    Number3[9][14] = 4'hC;
    Number3[10][14] = 4'hC;
    Number3[11][14] = 4'hC;
    Number3[12][14] = 4'hC;
    Number3[13][14] = 4'hC;
    Number3[14][14] = 4'hC;
    Number3[15][14] = 4'hC;
    Number3[16][14] = 4'hC;
    Number3[17][14] = 4'hD;
    Number3[18][14] = 4'hF;
    Number3[19][14] = 4'hF;
    Number3[20][14] = 4'hF;
    Number3[21][14] = 4'hF;
    Number3[22][14] = 4'hF;
    Number3[0][15] = 4'hF;
    Number3[1][15] = 4'hF;
    Number3[2][15] = 4'hF;
    Number3[3][15] = 4'hF;
    Number3[4][15] = 4'hF;
    Number3[5][15] = 4'hD;
    Number3[6][15] = 4'hC;
    Number3[7][15] = 4'hC;
    Number3[8][15] = 4'hC;
    Number3[9][15] = 4'hC;
    Number3[10][15] = 4'hC;
    Number3[11][15] = 4'hC;
    Number3[12][15] = 4'hC;
    Number3[13][15] = 4'hC;
    Number3[14][15] = 4'hC;
    Number3[15][15] = 4'hC;
    Number3[16][15] = 4'hC;
    Number3[17][15] = 4'hC;
    Number3[18][15] = 4'hD;
    Number3[19][15] = 4'hF;
    Number3[20][15] = 4'hF;
    Number3[21][15] = 4'hF;
    Number3[22][15] = 4'hF;
    Number3[0][16] = 4'hF;
    Number3[1][16] = 4'hF;
    Number3[2][16] = 4'hF;
    Number3[3][16] = 4'hF;
    Number3[4][16] = 4'hF;
    Number3[5][16] = 4'hF;
    Number3[6][16] = 4'hF;
    Number3[7][16] = 4'hF;
    Number3[8][16] = 4'hF;
    Number3[9][16] = 4'hF;
    Number3[10][16] = 4'hE;
    Number3[11][16] = 4'hD;
    Number3[12][16] = 4'hC;
    Number3[13][16] = 4'hC;
    Number3[14][16] = 4'hC;
    Number3[15][16] = 4'hC;
    Number3[16][16] = 4'hC;
    Number3[17][16] = 4'hC;
    Number3[18][16] = 4'hC;
    Number3[19][16] = 4'hD;
    Number3[20][16] = 4'hF;
    Number3[21][16] = 4'hF;
    Number3[22][16] = 4'hF;
    Number3[0][17] = 4'hF;
    Number3[1][17] = 4'hF;
    Number3[2][17] = 4'hF;
    Number3[3][17] = 4'hF;
    Number3[4][17] = 4'hF;
    Number3[5][17] = 4'hF;
    Number3[6][17] = 4'hF;
    Number3[7][17] = 4'hF;
    Number3[8][17] = 4'hF;
    Number3[9][17] = 4'hF;
    Number3[10][17] = 4'hF;
    Number3[11][17] = 4'hF;
    Number3[12][17] = 4'hF;
    Number3[13][17] = 4'hD;
    Number3[14][17] = 4'hC;
    Number3[15][17] = 4'hC;
    Number3[16][17] = 4'hC;
    Number3[17][17] = 4'hC;
    Number3[18][17] = 4'hC;
    Number3[19][17] = 4'hC;
    Number3[20][17] = 4'hF;
    Number3[21][17] = 4'hF;
    Number3[22][17] = 4'hF;
    Number3[0][18] = 4'hF;
    Number3[1][18] = 4'hF;
    Number3[2][18] = 4'hF;
    Number3[3][18] = 4'hF;
    Number3[4][18] = 4'hF;
    Number3[5][18] = 4'hF;
    Number3[6][18] = 4'hF;
    Number3[7][18] = 4'hF;
    Number3[8][18] = 4'hF;
    Number3[9][18] = 4'hF;
    Number3[10][18] = 4'hF;
    Number3[11][18] = 4'hF;
    Number3[12][18] = 4'hF;
    Number3[13][18] = 4'hE;
    Number3[14][18] = 4'hC;
    Number3[15][18] = 4'hC;
    Number3[16][18] = 4'hC;
    Number3[17][18] = 4'hC;
    Number3[18][18] = 4'hC;
    Number3[19][18] = 4'hC;
    Number3[20][18] = 4'hF;
    Number3[21][18] = 4'hF;
    Number3[22][18] = 4'hF;
    Number3[0][19] = 4'hF;
    Number3[1][19] = 4'hF;
    Number3[2][19] = 4'hF;
    Number3[3][19] = 4'hF;
    Number3[4][19] = 4'hF;
    Number3[5][19] = 4'hF;
    Number3[6][19] = 4'hF;
    Number3[7][19] = 4'hF;
    Number3[8][19] = 4'hF;
    Number3[9][19] = 4'hF;
    Number3[10][19] = 4'hF;
    Number3[11][19] = 4'hF;
    Number3[12][19] = 4'hF;
    Number3[13][19] = 4'hF;
    Number3[14][19] = 4'hC;
    Number3[15][19] = 4'hC;
    Number3[16][19] = 4'hC;
    Number3[17][19] = 4'hC;
    Number3[18][19] = 4'hC;
    Number3[19][19] = 4'hC;
    Number3[20][19] = 4'hF;
    Number3[21][19] = 4'hF;
    Number3[22][19] = 4'hF;
    Number3[0][20] = 4'hF;
    Number3[1][20] = 4'hF;
    Number3[2][20] = 4'hF;
    Number3[3][20] = 4'hF;
    Number3[4][20] = 4'hF;
    Number3[5][20] = 4'hF;
    Number3[6][20] = 4'hF;
    Number3[7][20] = 4'hF;
    Number3[8][20] = 4'hF;
    Number3[9][20] = 4'hF;
    Number3[10][20] = 4'hF;
    Number3[11][20] = 4'hF;
    Number3[12][20] = 4'hF;
    Number3[13][20] = 4'hF;
    Number3[14][20] = 4'hC;
    Number3[15][20] = 4'hC;
    Number3[16][20] = 4'hC;
    Number3[17][20] = 4'hC;
    Number3[18][20] = 4'hC;
    Number3[19][20] = 4'hC;
    Number3[20][20] = 4'hF;
    Number3[21][20] = 4'hF;
    Number3[22][20] = 4'hF;
    Number3[0][21] = 4'hF;
    Number3[1][21] = 4'hF;
    Number3[2][21] = 4'hF;
    Number3[3][21] = 4'hD;
    Number3[4][21] = 4'hD;
    Number3[5][21] = 4'hE;
    Number3[6][21] = 4'hF;
    Number3[7][21] = 4'hF;
    Number3[8][21] = 4'hF;
    Number3[9][21] = 4'hF;
    Number3[10][21] = 4'hF;
    Number3[11][21] = 4'hF;
    Number3[12][21] = 4'hF;
    Number3[13][21] = 4'hD;
    Number3[14][21] = 4'hC;
    Number3[15][21] = 4'hC;
    Number3[16][21] = 4'hC;
    Number3[17][21] = 4'hC;
    Number3[18][21] = 4'hC;
    Number3[19][21] = 4'hC;
    Number3[20][21] = 4'hF;
    Number3[21][21] = 4'hF;
    Number3[22][21] = 4'hF;
    Number3[0][22] = 4'hF;
    Number3[1][22] = 4'hF;
    Number3[2][22] = 4'hF;
    Number3[3][22] = 4'hC;
    Number3[4][22] = 4'hC;
    Number3[5][22] = 4'hC;
    Number3[6][22] = 4'hD;
    Number3[7][22] = 4'hD;
    Number3[8][22] = 4'hE;
    Number3[9][22] = 4'hF;
    Number3[10][22] = 4'hF;
    Number3[11][22] = 4'hE;
    Number3[12][22] = 4'hD;
    Number3[13][22] = 4'hC;
    Number3[14][22] = 4'hC;
    Number3[15][22] = 4'hC;
    Number3[16][22] = 4'hC;
    Number3[17][22] = 4'hC;
    Number3[18][22] = 4'hC;
    Number3[19][22] = 4'hD;
    Number3[20][22] = 4'hF;
    Number3[21][22] = 4'hF;
    Number3[22][22] = 4'hF;
    Number3[0][23] = 4'hF;
    Number3[1][23] = 4'hF;
    Number3[2][23] = 4'hF;
    Number3[3][23] = 4'hC;
    Number3[4][23] = 4'hC;
    Number3[5][23] = 4'hC;
    Number3[6][23] = 4'hC;
    Number3[7][23] = 4'hC;
    Number3[8][23] = 4'hC;
    Number3[9][23] = 4'hC;
    Number3[10][23] = 4'hC;
    Number3[11][23] = 4'hC;
    Number3[12][23] = 4'hC;
    Number3[13][23] = 4'hC;
    Number3[14][23] = 4'hC;
    Number3[15][23] = 4'hC;
    Number3[16][23] = 4'hC;
    Number3[17][23] = 4'hC;
    Number3[18][23] = 4'hC;
    Number3[19][23] = 4'hF;
    Number3[20][23] = 4'hF;
    Number3[21][23] = 4'hF;
    Number3[22][23] = 4'hF;
    Number3[0][24] = 4'hF;
    Number3[1][24] = 4'hF;
    Number3[2][24] = 4'hF;
    Number3[3][24] = 4'hD;
    Number3[4][24] = 4'hC;
    Number3[5][24] = 4'hC;
    Number3[6][24] = 4'hC;
    Number3[7][24] = 4'hC;
    Number3[8][24] = 4'hC;
    Number3[9][24] = 4'hC;
    Number3[10][24] = 4'hC;
    Number3[11][24] = 4'hC;
    Number3[12][24] = 4'hC;
    Number3[13][24] = 4'hC;
    Number3[14][24] = 4'hC;
    Number3[15][24] = 4'hC;
    Number3[16][24] = 4'hC;
    Number3[17][24] = 4'hC;
    Number3[18][24] = 4'hE;
    Number3[19][24] = 4'hF;
    Number3[20][24] = 4'hF;
    Number3[21][24] = 4'hF;
    Number3[22][24] = 4'hF;
    Number3[0][25] = 4'hF;
    Number3[1][25] = 4'hF;
    Number3[2][25] = 4'hF;
    Number3[3][25] = 4'hF;
    Number3[4][25] = 4'hD;
    Number3[5][25] = 4'hC;
    Number3[6][25] = 4'hC;
    Number3[7][25] = 4'hC;
    Number3[8][25] = 4'hC;
    Number3[9][25] = 4'hC;
    Number3[10][25] = 4'hC;
    Number3[11][25] = 4'hC;
    Number3[12][25] = 4'hC;
    Number3[13][25] = 4'hC;
    Number3[14][25] = 4'hC;
    Number3[15][25] = 4'hC;
    Number3[16][25] = 4'hD;
    Number3[17][25] = 4'hF;
    Number3[18][25] = 4'hF;
    Number3[19][25] = 4'hF;
    Number3[20][25] = 4'hF;
    Number3[21][25] = 4'hF;
    Number3[22][25] = 4'hF;
    Number3[0][26] = 4'hF;
    Number3[1][26] = 4'hF;
    Number3[2][26] = 4'hF;
    Number3[3][26] = 4'hF;
    Number3[4][26] = 4'hF;
    Number3[5][26] = 4'hF;
    Number3[6][26] = 4'hD;
    Number3[7][26] = 4'hD;
    Number3[8][26] = 4'hC;
    Number3[9][26] = 4'hC;
    Number3[10][26] = 4'hC;
    Number3[11][26] = 4'hC;
    Number3[12][26] = 4'hC;
    Number3[13][26] = 4'hD;
    Number3[14][26] = 4'hD;
    Number3[15][26] = 4'hE;
    Number3[16][26] = 4'hF;
    Number3[17][26] = 4'hF;
    Number3[18][26] = 4'hF;
    Number3[19][26] = 4'hF;
    Number3[20][26] = 4'hF;
    Number3[21][26] = 4'hF;
    Number3[22][26] = 4'hF;
    Number3[0][27] = 4'hF;
    Number3[1][27] = 4'hF;
    Number3[2][27] = 4'hF;
    Number3[3][27] = 4'hF;
    Number3[4][27] = 4'hF;
    Number3[5][27] = 4'hF;
    Number3[6][27] = 4'hF;
    Number3[7][27] = 4'hF;
    Number3[8][27] = 4'hF;
    Number3[9][27] = 4'hF;
    Number3[10][27] = 4'hF;
    Number3[11][27] = 4'hF;
    Number3[12][27] = 4'hF;
    Number3[13][27] = 4'hF;
    Number3[14][27] = 4'hF;
    Number3[15][27] = 4'hF;
    Number3[16][27] = 4'hF;
    Number3[17][27] = 4'hF;
    Number3[18][27] = 4'hF;
    Number3[19][27] = 4'hF;
    Number3[20][27] = 4'hF;
    Number3[21][27] = 4'hF;
    Number3[22][27] = 4'hF;
    Number3[0][28] = 4'hF;
    Number3[1][28] = 4'hF;
    Number3[2][28] = 4'hF;
    Number3[3][28] = 4'hF;
    Number3[4][28] = 4'hF;
    Number3[5][28] = 4'hF;
    Number3[6][28] = 4'hF;
    Number3[7][28] = 4'hF;
    Number3[8][28] = 4'hF;
    Number3[9][28] = 4'hF;
    Number3[10][28] = 4'hF;
    Number3[11][28] = 4'hF;
    Number3[12][28] = 4'hF;
    Number3[13][28] = 4'hF;
    Number3[14][28] = 4'hF;
    Number3[15][28] = 4'hF;
    Number3[16][28] = 4'hF;
    Number3[17][28] = 4'hF;
    Number3[18][28] = 4'hF;
    Number3[19][28] = 4'hF;
    Number3[20][28] = 4'hF;
    Number3[21][28] = 4'hF;
    Number3[22][28] = 4'hF;

// Number 4
    Number4[0][0] = 4'hF;
    Number4[1][0] = 4'hF;
    Number4[2][0] = 4'hF;
    Number4[3][0] = 4'hF;
    Number4[4][0] = 4'hF;
    Number4[5][0] = 4'hF;
    Number4[6][0] = 4'hF;
    Number4[7][0] = 4'hF;
    Number4[8][0] = 4'hF;
    Number4[9][0] = 4'hF;
    Number4[10][0] = 4'hF;
    Number4[11][0] = 4'hF;
    Number4[12][0] = 4'hF;
    Number4[13][0] = 4'hF;
    Number4[14][0] = 4'hF;
    Number4[15][0] = 4'hF;
    Number4[16][0] = 4'hF;
    Number4[17][0] = 4'hF;
    Number4[18][0] = 4'hF;
    Number4[19][0] = 4'hF;
    Number4[20][0] = 4'hF;
    Number4[21][0] = 4'hF;
    Number4[22][0] = 4'hF;
    Number4[0][1] = 4'hF;
    Number4[1][1] = 4'hF;
    Number4[2][1] = 4'hF;
    Number4[3][1] = 4'hF;
    Number4[4][1] = 4'hF;
    Number4[5][1] = 4'hF;
    Number4[6][1] = 4'hF;
    Number4[7][1] = 4'hF;
    Number4[8][1] = 4'hF;
    Number4[9][1] = 4'hF;
    Number4[10][1] = 4'hF;
    Number4[11][1] = 4'hF;
    Number4[12][1] = 4'hF;
    Number4[13][1] = 4'hF;
    Number4[14][1] = 4'hF;
    Number4[15][1] = 4'hF;
    Number4[16][1] = 4'hF;
    Number4[17][1] = 4'hF;
    Number4[18][1] = 4'hF;
    Number4[19][1] = 4'hF;
    Number4[20][1] = 4'hF;
    Number4[21][1] = 4'hF;
    Number4[22][1] = 4'hF;
    Number4[0][2] = 4'hF;
    Number4[1][2] = 4'hF;
    Number4[2][2] = 4'hF;
    Number4[3][2] = 4'hF;
    Number4[4][2] = 4'hF;
    Number4[5][2] = 4'hF;
    Number4[6][2] = 4'hF;
    Number4[7][2] = 4'hF;
    Number4[8][2] = 4'hF;
    Number4[9][2] = 4'hF;
    Number4[10][2] = 4'hE;
    Number4[11][2] = 4'hC;
    Number4[12][2] = 4'hC;
    Number4[13][2] = 4'hC;
    Number4[14][2] = 4'hC;
    Number4[15][2] = 4'hC;
    Number4[16][2] = 4'hC;
    Number4[17][2] = 4'hD;
    Number4[18][2] = 4'hF;
    Number4[19][2] = 4'hF;
    Number4[20][2] = 4'hF;
    Number4[21][2] = 4'hF;
    Number4[22][2] = 4'hF;
    Number4[0][3] = 4'hF;
    Number4[1][3] = 4'hF;
    Number4[2][3] = 4'hF;
    Number4[3][3] = 4'hF;
    Number4[4][3] = 4'hF;
    Number4[5][3] = 4'hF;
    Number4[6][3] = 4'hF;
    Number4[7][3] = 4'hF;
    Number4[8][3] = 4'hF;
    Number4[9][3] = 4'hF;
    Number4[10][3] = 4'hC;
    Number4[11][3] = 4'hC;
    Number4[12][3] = 4'hC;
    Number4[13][3] = 4'hC;
    Number4[14][3] = 4'hC;
    Number4[15][3] = 4'hC;
    Number4[16][3] = 4'hC;
    Number4[17][3] = 4'hC;
    Number4[18][3] = 4'hF;
    Number4[19][3] = 4'hF;
    Number4[20][3] = 4'hF;
    Number4[21][3] = 4'hF;
    Number4[22][3] = 4'hF;
    Number4[0][4] = 4'hF;
    Number4[1][4] = 4'hF;
    Number4[2][4] = 4'hF;
    Number4[3][4] = 4'hF;
    Number4[4][4] = 4'hF;
    Number4[5][4] = 4'hF;
    Number4[6][4] = 4'hF;
    Number4[7][4] = 4'hF;
    Number4[8][4] = 4'hF;
    Number4[9][4] = 4'hD;
    Number4[10][4] = 4'hC;
    Number4[11][4] = 4'hC;
    Number4[12][4] = 4'hC;
    Number4[13][4] = 4'hC;
    Number4[14][4] = 4'hC;
    Number4[15][4] = 4'hC;
    Number4[16][4] = 4'hC;
    Number4[17][4] = 4'hC;
    Number4[18][4] = 4'hF;
    Number4[19][4] = 4'hF;
    Number4[20][4] = 4'hF;
    Number4[21][4] = 4'hF;
    Number4[22][4] = 4'hF;
    Number4[0][5] = 4'hF;
    Number4[1][5] = 4'hF;
    Number4[2][5] = 4'hF;
    Number4[3][5] = 4'hF;
    Number4[4][5] = 4'hF;
    Number4[5][5] = 4'hF;
    Number4[6][5] = 4'hF;
    Number4[7][5] = 4'hF;
    Number4[8][5] = 4'hF;
    Number4[9][5] = 4'hC;
    Number4[10][5] = 4'hC;
    Number4[11][5] = 4'hC;
    Number4[12][5] = 4'hC;
    Number4[13][5] = 4'hC;
    Number4[14][5] = 4'hC;
    Number4[15][5] = 4'hC;
    Number4[16][5] = 4'hC;
    Number4[17][5] = 4'hC;
    Number4[18][5] = 4'hF;
    Number4[19][5] = 4'hF;
    Number4[20][5] = 4'hF;
    Number4[21][5] = 4'hF;
    Number4[22][5] = 4'hF;
    Number4[0][6] = 4'hF;
    Number4[1][6] = 4'hF;
    Number4[2][6] = 4'hF;
    Number4[3][6] = 4'hF;
    Number4[4][6] = 4'hF;
    Number4[5][6] = 4'hF;
    Number4[6][6] = 4'hF;
    Number4[7][6] = 4'hF;
    Number4[8][6] = 4'hD;
    Number4[9][6] = 4'hC;
    Number4[10][6] = 4'hC;
    Number4[11][6] = 4'hC;
    Number4[12][6] = 4'hD;
    Number4[13][6] = 4'hC;
    Number4[14][6] = 4'hC;
    Number4[15][6] = 4'hC;
    Number4[16][6] = 4'hC;
    Number4[17][6] = 4'hC;
    Number4[18][6] = 4'hF;
    Number4[19][6] = 4'hF;
    Number4[20][6] = 4'hF;
    Number4[21][6] = 4'hF;
    Number4[22][6] = 4'hF;
    Number4[0][7] = 4'hF;
    Number4[1][7] = 4'hF;
    Number4[2][7] = 4'hF;
    Number4[3][7] = 4'hF;
    Number4[4][7] = 4'hF;
    Number4[5][7] = 4'hF;
    Number4[6][7] = 4'hF;
    Number4[7][7] = 4'hE;
    Number4[8][7] = 4'hC;
    Number4[9][7] = 4'hC;
    Number4[10][7] = 4'hC;
    Number4[11][7] = 4'hC;
    Number4[12][7] = 4'hE;
    Number4[13][7] = 4'hC;
    Number4[14][7] = 4'hC;
    Number4[15][7] = 4'hC;
    Number4[16][7] = 4'hC;
    Number4[17][7] = 4'hC;
    Number4[18][7] = 4'hF;
    Number4[19][7] = 4'hF;
    Number4[20][7] = 4'hF;
    Number4[21][7] = 4'hF;
    Number4[22][7] = 4'hF;
    Number4[0][8] = 4'hF;
    Number4[1][8] = 4'hF;
    Number4[2][8] = 4'hF;
    Number4[3][8] = 4'hF;
    Number4[4][8] = 4'hF;
    Number4[5][8] = 4'hF;
    Number4[6][8] = 4'hF;
    Number4[7][8] = 4'hD;
    Number4[8][8] = 4'hC;
    Number4[9][8] = 4'hC;
    Number4[10][8] = 4'hC;
    Number4[11][8] = 4'hD;
    Number4[12][8] = 4'hF;
    Number4[13][8] = 4'hC;
    Number4[14][8] = 4'hC;
    Number4[15][8] = 4'hC;
    Number4[16][8] = 4'hC;
    Number4[17][8] = 4'hC;
    Number4[18][8] = 4'hF;
    Number4[19][8] = 4'hF;
    Number4[20][8] = 4'hF;
    Number4[21][8] = 4'hF;
    Number4[22][8] = 4'hF;
    Number4[0][9] = 4'hF;
    Number4[1][9] = 4'hF;
    Number4[2][9] = 4'hF;
    Number4[3][9] = 4'hF;
    Number4[4][9] = 4'hF;
    Number4[5][9] = 4'hF;
    Number4[6][9] = 4'hE;
    Number4[7][9] = 4'hC;
    Number4[8][9] = 4'hC;
    Number4[9][9] = 4'hC;
    Number4[10][9] = 4'hC;
    Number4[11][9] = 4'hE;
    Number4[12][9] = 4'hF;
    Number4[13][9] = 4'hC;
    Number4[14][9] = 4'hC;
    Number4[15][9] = 4'hC;
    Number4[16][9] = 4'hC;
    Number4[17][9] = 4'hC;
    Number4[18][9] = 4'hF;
    Number4[19][9] = 4'hF;
    Number4[20][9] = 4'hF;
    Number4[21][9] = 4'hF;
    Number4[22][9] = 4'hF;
    Number4[0][10] = 4'hF;
    Number4[1][10] = 4'hF;
    Number4[2][10] = 4'hF;
    Number4[3][10] = 4'hF;
    Number4[4][10] = 4'hF;
    Number4[5][10] = 4'hF;
    Number4[6][10] = 4'hC;
    Number4[7][10] = 4'hC;
    Number4[8][10] = 4'hC;
    Number4[9][10] = 4'hC;
    Number4[10][10] = 4'hD;
    Number4[11][10] = 4'hF;
    Number4[12][10] = 4'hF;
    Number4[13][10] = 4'hC;
    Number4[14][10] = 4'hC;
    Number4[15][10] = 4'hC;
    Number4[16][10] = 4'hC;
    Number4[17][10] = 4'hC;
    Number4[18][10] = 4'hF;
    Number4[19][10] = 4'hF;
    Number4[20][10] = 4'hF;
    Number4[21][10] = 4'hF;
    Number4[22][10] = 4'hF;
    Number4[0][11] = 4'hF;
    Number4[1][11] = 4'hF;
    Number4[2][11] = 4'hF;
    Number4[3][11] = 4'hF;
    Number4[4][11] = 4'hF;
    Number4[5][11] = 4'hD;
    Number4[6][11] = 4'hC;
    Number4[7][11] = 4'hC;
    Number4[8][11] = 4'hC;
    Number4[9][11] = 4'hC;
    Number4[10][11] = 4'hF;
    Number4[11][11] = 4'hF;
    Number4[12][11] = 4'hF;
    Number4[13][11] = 4'hC;
    Number4[14][11] = 4'hC;
    Number4[15][11] = 4'hC;
    Number4[16][11] = 4'hC;
    Number4[17][11] = 4'hC;
    Number4[18][11] = 4'hF;
    Number4[19][11] = 4'hF;
    Number4[20][11] = 4'hF;
    Number4[21][11] = 4'hF;
    Number4[22][11] = 4'hF;
    Number4[0][12] = 4'hF;
    Number4[1][12] = 4'hF;
    Number4[2][12] = 4'hF;
    Number4[3][12] = 4'hF;
    Number4[4][12] = 4'hF;
    Number4[5][12] = 4'hC;
    Number4[6][12] = 4'hC;
    Number4[7][12] = 4'hC;
    Number4[8][12] = 4'hC;
    Number4[9][12] = 4'hD;
    Number4[10][12] = 4'hF;
    Number4[11][12] = 4'hF;
    Number4[12][12] = 4'hF;
    Number4[13][12] = 4'hC;
    Number4[14][12] = 4'hC;
    Number4[15][12] = 4'hC;
    Number4[16][12] = 4'hC;
    Number4[17][12] = 4'hC;
    Number4[18][12] = 4'hF;
    Number4[19][12] = 4'hF;
    Number4[20][12] = 4'hF;
    Number4[21][12] = 4'hF;
    Number4[22][12] = 4'hF;
    Number4[0][13] = 4'hF;
    Number4[1][13] = 4'hF;
    Number4[2][13] = 4'hF;
    Number4[3][13] = 4'hF;
    Number4[4][13] = 4'hD;
    Number4[5][13] = 4'hC;
    Number4[6][13] = 4'hC;
    Number4[7][13] = 4'hC;
    Number4[8][13] = 4'hC;
    Number4[9][13] = 4'hF;
    Number4[10][13] = 4'hF;
    Number4[11][13] = 4'hF;
    Number4[12][13] = 4'hF;
    Number4[13][13] = 4'hC;
    Number4[14][13] = 4'hC;
    Number4[15][13] = 4'hC;
    Number4[16][13] = 4'hC;
    Number4[17][13] = 4'hC;
    Number4[18][13] = 4'hF;
    Number4[19][13] = 4'hF;
    Number4[20][13] = 4'hF;
    Number4[21][13] = 4'hF;
    Number4[22][13] = 4'hF;
    Number4[0][14] = 4'hF;
    Number4[1][14] = 4'hF;
    Number4[2][14] = 4'hF;
    Number4[3][14] = 4'hE;
    Number4[4][14] = 4'hC;
    Number4[5][14] = 4'hC;
    Number4[6][14] = 4'hC;
    Number4[7][14] = 4'hC;
    Number4[8][14] = 4'hD;
    Number4[9][14] = 4'hF;
    Number4[10][14] = 4'hF;
    Number4[11][14] = 4'hF;
    Number4[12][14] = 4'hF;
    Number4[13][14] = 4'hC;
    Number4[14][14] = 4'hC;
    Number4[15][14] = 4'hC;
    Number4[16][14] = 4'hC;
    Number4[17][14] = 4'hC;
    Number4[18][14] = 4'hF;
    Number4[19][14] = 4'hF;
    Number4[20][14] = 4'hF;
    Number4[21][14] = 4'hF;
    Number4[22][14] = 4'hF;
    Number4[0][15] = 4'hF;
    Number4[1][15] = 4'hF;
    Number4[2][15] = 4'hF;
    Number4[3][15] = 4'hD;
    Number4[4][15] = 4'hC;
    Number4[5][15] = 4'hC;
    Number4[6][15] = 4'hC;
    Number4[7][15] = 4'hC;
    Number4[8][15] = 4'hF;
    Number4[9][15] = 4'hF;
    Number4[10][15] = 4'hF;
    Number4[11][15] = 4'hF;
    Number4[12][15] = 4'hF;
    Number4[13][15] = 4'hC;
    Number4[14][15] = 4'hC;
    Number4[15][15] = 4'hC;
    Number4[16][15] = 4'hC;
    Number4[17][15] = 4'hC;
    Number4[18][15] = 4'hF;
    Number4[19][15] = 4'hF;
    Number4[20][15] = 4'hF;
    Number4[21][15] = 4'hF;
    Number4[22][15] = 4'hF;
    Number4[0][16] = 4'hF;
    Number4[1][16] = 4'hF;
    Number4[2][16] = 4'hE;
    Number4[3][16] = 4'hC;
    Number4[4][16] = 4'hC;
    Number4[5][16] = 4'hC;
    Number4[6][16] = 4'hC;
    Number4[7][16] = 4'hE;
    Number4[8][16] = 4'hF;
    Number4[9][16] = 4'hF;
    Number4[10][16] = 4'hF;
    Number4[11][16] = 4'hF;
    Number4[12][16] = 4'hF;
    Number4[13][16] = 4'hC;
    Number4[14][16] = 4'hC;
    Number4[15][16] = 4'hC;
    Number4[16][16] = 4'hC;
    Number4[17][16] = 4'hC;
    Number4[18][16] = 4'hF;
    Number4[19][16] = 4'hF;
    Number4[20][16] = 4'hF;
    Number4[21][16] = 4'hF;
    Number4[22][16] = 4'hF;
    Number4[0][17] = 4'hF;
    Number4[1][17] = 4'hF;
    Number4[2][17] = 4'hD;
    Number4[3][17] = 4'hC;
    Number4[4][17] = 4'hC;
    Number4[5][17] = 4'hC;
    Number4[6][17] = 4'hD;
    Number4[7][17] = 4'hF;
    Number4[8][17] = 4'hF;
    Number4[9][17] = 4'hF;
    Number4[10][17] = 4'hF;
    Number4[11][17] = 4'hF;
    Number4[12][17] = 4'hF;
    Number4[13][17] = 4'hC;
    Number4[14][17] = 4'hC;
    Number4[15][17] = 4'hC;
    Number4[16][17] = 4'hC;
    Number4[17][17] = 4'hC;
    Number4[18][17] = 4'hF;
    Number4[19][17] = 4'hF;
    Number4[20][17] = 4'hF;
    Number4[21][17] = 4'hF;
    Number4[22][17] = 4'hF;
    Number4[0][18] = 4'hF;
    Number4[1][18] = 4'hF;
    Number4[2][18] = 4'hC;
    Number4[3][18] = 4'hC;
    Number4[4][18] = 4'hC;
    Number4[5][18] = 4'hC;
    Number4[6][18] = 4'hC;
    Number4[7][18] = 4'hC;
    Number4[8][18] = 4'hC;
    Number4[9][18] = 4'hC;
    Number4[10][18] = 4'hC;
    Number4[11][18] = 4'hC;
    Number4[12][18] = 4'hC;
    Number4[13][18] = 4'hC;
    Number4[14][18] = 4'hC;
    Number4[15][18] = 4'hC;
    Number4[16][18] = 4'hC;
    Number4[17][18] = 4'hC;
    Number4[18][18] = 4'hC;
    Number4[19][18] = 4'hC;
    Number4[20][18] = 4'hD;
    Number4[21][18] = 4'hF;
    Number4[22][18] = 4'hF;
    Number4[0][19] = 4'hF;
    Number4[1][19] = 4'hF;
    Number4[2][19] = 4'hC;
    Number4[3][19] = 4'hC;
    Number4[4][19] = 4'hC;
    Number4[5][19] = 4'hC;
    Number4[6][19] = 4'hC;
    Number4[7][19] = 4'hC;
    Number4[8][19] = 4'hC;
    Number4[9][19] = 4'hC;
    Number4[10][19] = 4'hC;
    Number4[11][19] = 4'hC;
    Number4[12][19] = 4'hC;
    Number4[13][19] = 4'hC;
    Number4[14][19] = 4'hC;
    Number4[15][19] = 4'hC;
    Number4[16][19] = 4'hC;
    Number4[17][19] = 4'hC;
    Number4[18][19] = 4'hC;
    Number4[19][19] = 4'hC;
    Number4[20][19] = 4'hC;
    Number4[21][19] = 4'hF;
    Number4[22][19] = 4'hF;
    Number4[0][20] = 4'hF;
    Number4[1][20] = 4'hF;
    Number4[2][20] = 4'hC;
    Number4[3][20] = 4'hC;
    Number4[4][20] = 4'hC;
    Number4[5][20] = 4'hC;
    Number4[6][20] = 4'hC;
    Number4[7][20] = 4'hC;
    Number4[8][20] = 4'hC;
    Number4[9][20] = 4'hC;
    Number4[10][20] = 4'hC;
    Number4[11][20] = 4'hC;
    Number4[12][20] = 4'hC;
    Number4[13][20] = 4'hC;
    Number4[14][20] = 4'hC;
    Number4[15][20] = 4'hC;
    Number4[16][20] = 4'hC;
    Number4[17][20] = 4'hC;
    Number4[18][20] = 4'hC;
    Number4[19][20] = 4'hC;
    Number4[20][20] = 4'hC;
    Number4[21][20] = 4'hF;
    Number4[22][20] = 4'hF;
    Number4[0][21] = 4'hF;
    Number4[1][21] = 4'hF;
    Number4[2][21] = 4'hD;
    Number4[3][21] = 4'hC;
    Number4[4][21] = 4'hC;
    Number4[5][21] = 4'hC;
    Number4[6][21] = 4'hC;
    Number4[7][21] = 4'hC;
    Number4[8][21] = 4'hC;
    Number4[9][21] = 4'hC;
    Number4[10][21] = 4'hC;
    Number4[11][21] = 4'hC;
    Number4[12][21] = 4'hC;
    Number4[13][21] = 4'hC;
    Number4[14][21] = 4'hC;
    Number4[15][21] = 4'hC;
    Number4[16][21] = 4'hC;
    Number4[17][21] = 4'hC;
    Number4[18][21] = 4'hC;
    Number4[19][21] = 4'hC;
    Number4[20][21] = 4'hD;
    Number4[21][21] = 4'hF;
    Number4[22][21] = 4'hF;
    Number4[0][22] = 4'hF;
    Number4[1][22] = 4'hF;
    Number4[2][22] = 4'hF;
    Number4[3][22] = 4'hF;
    Number4[4][22] = 4'hF;
    Number4[5][22] = 4'hF;
    Number4[6][22] = 4'hF;
    Number4[7][22] = 4'hF;
    Number4[8][22] = 4'hF;
    Number4[9][22] = 4'hF;
    Number4[10][22] = 4'hF;
    Number4[11][22] = 4'hF;
    Number4[12][22] = 4'hF;
    Number4[13][22] = 4'hC;
    Number4[14][22] = 4'hC;
    Number4[15][22] = 4'hC;
    Number4[16][22] = 4'hC;
    Number4[17][22] = 4'hC;
    Number4[18][22] = 4'hF;
    Number4[19][22] = 4'hF;
    Number4[20][22] = 4'hF;
    Number4[21][22] = 4'hF;
    Number4[22][22] = 4'hF;
    Number4[0][23] = 4'hF;
    Number4[1][23] = 4'hF;
    Number4[2][23] = 4'hF;
    Number4[3][23] = 4'hF;
    Number4[4][23] = 4'hF;
    Number4[5][23] = 4'hF;
    Number4[6][23] = 4'hF;
    Number4[7][23] = 4'hF;
    Number4[8][23] = 4'hF;
    Number4[9][23] = 4'hF;
    Number4[10][23] = 4'hF;
    Number4[11][23] = 4'hF;
    Number4[12][23] = 4'hF;
    Number4[13][23] = 4'hC;
    Number4[14][23] = 4'hC;
    Number4[15][23] = 4'hC;
    Number4[16][23] = 4'hC;
    Number4[17][23] = 4'hC;
    Number4[18][23] = 4'hF;
    Number4[19][23] = 4'hF;
    Number4[20][23] = 4'hF;
    Number4[21][23] = 4'hF;
    Number4[22][23] = 4'hF;
    Number4[0][24] = 4'hF;
    Number4[1][24] = 4'hF;
    Number4[2][24] = 4'hF;
    Number4[3][24] = 4'hF;
    Number4[4][24] = 4'hF;
    Number4[5][24] = 4'hF;
    Number4[6][24] = 4'hF;
    Number4[7][24] = 4'hF;
    Number4[8][24] = 4'hF;
    Number4[9][24] = 4'hF;
    Number4[10][24] = 4'hF;
    Number4[11][24] = 4'hF;
    Number4[12][24] = 4'hF;
    Number4[13][24] = 4'hC;
    Number4[14][24] = 4'hC;
    Number4[15][24] = 4'hC;
    Number4[16][24] = 4'hC;
    Number4[17][24] = 4'hC;
    Number4[18][24] = 4'hF;
    Number4[19][24] = 4'hF;
    Number4[20][24] = 4'hF;
    Number4[21][24] = 4'hF;
    Number4[22][24] = 4'hF;
    Number4[0][25] = 4'hF;
    Number4[1][25] = 4'hF;
    Number4[2][25] = 4'hF;
    Number4[3][25] = 4'hF;
    Number4[4][25] = 4'hF;
    Number4[5][25] = 4'hF;
    Number4[6][25] = 4'hF;
    Number4[7][25] = 4'hF;
    Number4[8][25] = 4'hF;
    Number4[9][25] = 4'hF;
    Number4[10][25] = 4'hF;
    Number4[11][25] = 4'hF;
    Number4[12][25] = 4'hF;
    Number4[13][25] = 4'hC;
    Number4[14][25] = 4'hC;
    Number4[15][25] = 4'hC;
    Number4[16][25] = 4'hC;
    Number4[17][25] = 4'hC;
    Number4[18][25] = 4'hF;
    Number4[19][25] = 4'hF;
    Number4[20][25] = 4'hF;
    Number4[21][25] = 4'hF;
    Number4[22][25] = 4'hF;
    Number4[0][26] = 4'hF;
    Number4[1][26] = 4'hF;
    Number4[2][26] = 4'hF;
    Number4[3][26] = 4'hF;
    Number4[4][26] = 4'hF;
    Number4[5][26] = 4'hF;
    Number4[6][26] = 4'hF;
    Number4[7][26] = 4'hF;
    Number4[8][26] = 4'hF;
    Number4[9][26] = 4'hF;
    Number4[10][26] = 4'hF;
    Number4[11][26] = 4'hF;
    Number4[12][26] = 4'hF;
    Number4[13][26] = 4'hC;
    Number4[14][26] = 4'hC;
    Number4[15][26] = 4'hC;
    Number4[16][26] = 4'hC;
    Number4[17][26] = 4'hC;
    Number4[18][26] = 4'hF;
    Number4[19][26] = 4'hF;
    Number4[20][26] = 4'hF;
    Number4[21][26] = 4'hF;
    Number4[22][26] = 4'hF;
    Number4[0][27] = 4'hF;
    Number4[1][27] = 4'hF;
    Number4[2][27] = 4'hF;
    Number4[3][27] = 4'hF;
    Number4[4][27] = 4'hF;
    Number4[5][27] = 4'hF;
    Number4[6][27] = 4'hF;
    Number4[7][27] = 4'hF;
    Number4[8][27] = 4'hF;
    Number4[9][27] = 4'hF;
    Number4[10][27] = 4'hF;
    Number4[11][27] = 4'hF;
    Number4[12][27] = 4'hF;
    Number4[13][27] = 4'hF;
    Number4[14][27] = 4'hF;
    Number4[15][27] = 4'hF;
    Number4[16][27] = 4'hF;
    Number4[17][27] = 4'hF;
    Number4[18][27] = 4'hF;
    Number4[19][27] = 4'hF;
    Number4[20][27] = 4'hF;
    Number4[21][27] = 4'hF;
    Number4[22][27] = 4'hF;
    Number4[0][28] = 4'hF;
    Number4[1][28] = 4'hF;
    Number4[2][28] = 4'hF;
    Number4[3][28] = 4'hF;
    Number4[4][28] = 4'hF;
    Number4[5][28] = 4'hF;
    Number4[6][28] = 4'hF;
    Number4[7][28] = 4'hF;
    Number4[8][28] = 4'hF;
    Number4[9][28] = 4'hF;
    Number4[10][28] = 4'hF;
    Number4[11][28] = 4'hF;
    Number4[12][28] = 4'hF;
    Number4[13][28] = 4'hF;
    Number4[14][28] = 4'hF;
    Number4[15][28] = 4'hF;
    Number4[16][28] = 4'hF;
    Number4[17][28] = 4'hF;
    Number4[18][28] = 4'hF;
    Number4[19][28] = 4'hF;
    Number4[20][28] = 4'hF;
    Number4[21][28] = 4'hF;
    Number4[22][28] = 4'hF;

// Number 5
    Number5[0][0] = 4'hF;
    Number5[1][0] = 4'hF;
    Number5[2][0] = 4'hF;
    Number5[3][0] = 4'hF;
    Number5[4][0] = 4'hF;
    Number5[5][0] = 4'hF;
    Number5[6][0] = 4'hF;
    Number5[7][0] = 4'hF;
    Number5[8][0] = 4'hF;
    Number5[9][0] = 4'hF;
    Number5[10][0] = 4'hF;
    Number5[11][0] = 4'hF;
    Number5[12][0] = 4'hF;
    Number5[13][0] = 4'hF;
    Number5[14][0] = 4'hF;
    Number5[15][0] = 4'hF;
    Number5[16][0] = 4'hF;
    Number5[17][0] = 4'hF;
    Number5[18][0] = 4'hF;
    Number5[19][0] = 4'hF;
    Number5[20][0] = 4'hF;
    Number5[21][0] = 4'hF;
    Number5[22][0] = 4'hF;
    Number5[0][1] = 4'hF;
    Number5[1][1] = 4'hF;
    Number5[2][1] = 4'hF;
    Number5[3][1] = 4'hF;
    Number5[4][1] = 4'hF;
    Number5[5][1] = 4'hF;
    Number5[6][1] = 4'hF;
    Number5[7][1] = 4'hF;
    Number5[8][1] = 4'hF;
    Number5[9][1] = 4'hF;
    Number5[10][1] = 4'hF;
    Number5[11][1] = 4'hF;
    Number5[12][1] = 4'hF;
    Number5[13][1] = 4'hF;
    Number5[14][1] = 4'hF;
    Number5[15][1] = 4'hF;
    Number5[16][1] = 4'hF;
    Number5[17][1] = 4'hF;
    Number5[18][1] = 4'hF;
    Number5[19][1] = 4'hF;
    Number5[20][1] = 4'hF;
    Number5[21][1] = 4'hF;
    Number5[22][1] = 4'hF;
    Number5[0][2] = 4'hF;
    Number5[1][2] = 4'hF;
    Number5[2][2] = 4'hF;
    Number5[3][2] = 4'hF;
    Number5[4][2] = 4'hD;
    Number5[5][2] = 4'hC;
    Number5[6][2] = 4'hC;
    Number5[7][2] = 4'hC;
    Number5[8][2] = 4'hC;
    Number5[9][2] = 4'hC;
    Number5[10][2] = 4'hC;
    Number5[11][2] = 4'hC;
    Number5[12][2] = 4'hC;
    Number5[13][2] = 4'hC;
    Number5[14][2] = 4'hC;
    Number5[15][2] = 4'hC;
    Number5[16][2] = 4'hC;
    Number5[17][2] = 4'hC;
    Number5[18][2] = 4'hE;
    Number5[19][2] = 4'hF;
    Number5[20][2] = 4'hF;
    Number5[21][2] = 4'hF;
    Number5[22][2] = 4'hF;
    Number5[0][3] = 4'hF;
    Number5[1][3] = 4'hF;
    Number5[2][3] = 4'hF;
    Number5[3][3] = 4'hF;
    Number5[4][3] = 4'hD;
    Number5[5][3] = 4'hC;
    Number5[6][3] = 4'hC;
    Number5[7][3] = 4'hC;
    Number5[8][3] = 4'hC;
    Number5[9][3] = 4'hC;
    Number5[10][3] = 4'hC;
    Number5[11][3] = 4'hC;
    Number5[12][3] = 4'hC;
    Number5[13][3] = 4'hC;
    Number5[14][3] = 4'hC;
    Number5[15][3] = 4'hC;
    Number5[16][3] = 4'hC;
    Number5[17][3] = 4'hC;
    Number5[18][3] = 4'hD;
    Number5[19][3] = 4'hF;
    Number5[20][3] = 4'hF;
    Number5[21][3] = 4'hF;
    Number5[22][3] = 4'hF;
    Number5[0][4] = 4'hF;
    Number5[1][4] = 4'hF;
    Number5[2][4] = 4'hF;
    Number5[3][4] = 4'hF;
    Number5[4][4] = 4'hD;
    Number5[5][4] = 4'hC;
    Number5[6][4] = 4'hC;
    Number5[7][4] = 4'hC;
    Number5[8][4] = 4'hC;
    Number5[9][4] = 4'hC;
    Number5[10][4] = 4'hC;
    Number5[11][4] = 4'hC;
    Number5[12][4] = 4'hC;
    Number5[13][4] = 4'hC;
    Number5[14][4] = 4'hC;
    Number5[15][4] = 4'hC;
    Number5[16][4] = 4'hC;
    Number5[17][4] = 4'hC;
    Number5[18][4] = 4'hD;
    Number5[19][4] = 4'hF;
    Number5[20][4] = 4'hF;
    Number5[21][4] = 4'hF;
    Number5[22][4] = 4'hF;
    Number5[0][5] = 4'hF;
    Number5[1][5] = 4'hF;
    Number5[2][5] = 4'hF;
    Number5[3][5] = 4'hF;
    Number5[4][5] = 4'hD;
    Number5[5][5] = 4'hC;
    Number5[6][5] = 4'hC;
    Number5[7][5] = 4'hC;
    Number5[8][5] = 4'hC;
    Number5[9][5] = 4'hC;
    Number5[10][5] = 4'hC;
    Number5[11][5] = 4'hC;
    Number5[12][5] = 4'hC;
    Number5[13][5] = 4'hC;
    Number5[14][5] = 4'hC;
    Number5[15][5] = 4'hC;
    Number5[16][5] = 4'hC;
    Number5[17][5] = 4'hC;
    Number5[18][5] = 4'hE;
    Number5[19][5] = 4'hF;
    Number5[20][5] = 4'hF;
    Number5[21][5] = 4'hF;
    Number5[22][5] = 4'hF;
    Number5[0][6] = 4'hF;
    Number5[1][6] = 4'hF;
    Number5[2][6] = 4'hF;
    Number5[3][6] = 4'hF;
    Number5[4][6] = 4'hD;
    Number5[5][6] = 4'hC;
    Number5[6][6] = 4'hC;
    Number5[7][6] = 4'hC;
    Number5[8][6] = 4'hD;
    Number5[9][6] = 4'hF;
    Number5[10][6] = 4'hF;
    Number5[11][6] = 4'hF;
    Number5[12][6] = 4'hF;
    Number5[13][6] = 4'hF;
    Number5[14][6] = 4'hF;
    Number5[15][6] = 4'hF;
    Number5[16][6] = 4'hF;
    Number5[17][6] = 4'hF;
    Number5[18][6] = 4'hF;
    Number5[19][6] = 4'hF;
    Number5[20][6] = 4'hF;
    Number5[21][6] = 4'hF;
    Number5[22][6] = 4'hF;
    Number5[0][7] = 4'hF;
    Number5[1][7] = 4'hF;
    Number5[2][7] = 4'hF;
    Number5[3][7] = 4'hF;
    Number5[4][7] = 4'hD;
    Number5[5][7] = 4'hC;
    Number5[6][7] = 4'hC;
    Number5[7][7] = 4'hC;
    Number5[8][7] = 4'hD;
    Number5[9][7] = 4'hF;
    Number5[10][7] = 4'hF;
    Number5[11][7] = 4'hF;
    Number5[12][7] = 4'hF;
    Number5[13][7] = 4'hF;
    Number5[14][7] = 4'hF;
    Number5[15][7] = 4'hF;
    Number5[16][7] = 4'hF;
    Number5[17][7] = 4'hF;
    Number5[18][7] = 4'hF;
    Number5[19][7] = 4'hF;
    Number5[20][7] = 4'hF;
    Number5[21][7] = 4'hF;
    Number5[22][7] = 4'hF;
    Number5[0][8] = 4'hF;
    Number5[1][8] = 4'hF;
    Number5[2][8] = 4'hF;
    Number5[3][8] = 4'hF;
    Number5[4][8] = 4'hD;
    Number5[5][8] = 4'hC;
    Number5[6][8] = 4'hC;
    Number5[7][8] = 4'hC;
    Number5[8][8] = 4'hD;
    Number5[9][8] = 4'hF;
    Number5[10][8] = 4'hF;
    Number5[11][8] = 4'hF;
    Number5[12][8] = 4'hF;
    Number5[13][8] = 4'hF;
    Number5[14][8] = 4'hF;
    Number5[15][8] = 4'hF;
    Number5[16][8] = 4'hF;
    Number5[17][8] = 4'hF;
    Number5[18][8] = 4'hF;
    Number5[19][8] = 4'hF;
    Number5[20][8] = 4'hF;
    Number5[21][8] = 4'hF;
    Number5[22][8] = 4'hF;
    Number5[0][9] = 4'hF;
    Number5[1][9] = 4'hF;
    Number5[2][9] = 4'hF;
    Number5[3][9] = 4'hF;
    Number5[4][9] = 4'hD;
    Number5[5][9] = 4'hC;
    Number5[6][9] = 4'hC;
    Number5[7][9] = 4'hC;
    Number5[8][9] = 4'hD;
    Number5[9][9] = 4'hF;
    Number5[10][9] = 4'hF;
    Number5[11][9] = 4'hF;
    Number5[12][9] = 4'hF;
    Number5[13][9] = 4'hF;
    Number5[14][9] = 4'hF;
    Number5[15][9] = 4'hF;
    Number5[16][9] = 4'hF;
    Number5[17][9] = 4'hF;
    Number5[18][9] = 4'hF;
    Number5[19][9] = 4'hF;
    Number5[20][9] = 4'hF;
    Number5[21][9] = 4'hF;
    Number5[22][9] = 4'hF;
    Number5[0][10] = 4'hF;
    Number5[1][10] = 4'hF;
    Number5[2][10] = 4'hF;
    Number5[3][10] = 4'hF;
    Number5[4][10] = 4'hD;
    Number5[5][10] = 4'hC;
    Number5[6][10] = 4'hC;
    Number5[7][10] = 4'hC;
    Number5[8][10] = 4'hD;
    Number5[9][10] = 4'hF;
    Number5[10][10] = 4'hF;
    Number5[11][10] = 4'hF;
    Number5[12][10] = 4'hF;
    Number5[13][10] = 4'hF;
    Number5[14][10] = 4'hF;
    Number5[15][10] = 4'hF;
    Number5[16][10] = 4'hF;
    Number5[17][10] = 4'hF;
    Number5[18][10] = 4'hF;
    Number5[19][10] = 4'hF;
    Number5[20][10] = 4'hF;
    Number5[21][10] = 4'hF;
    Number5[22][10] = 4'hF;
    Number5[0][11] = 4'hF;
    Number5[1][11] = 4'hF;
    Number5[2][11] = 4'hF;
    Number5[3][11] = 4'hF;
    Number5[4][11] = 4'hD;
    Number5[5][11] = 4'hC;
    Number5[6][11] = 4'hC;
    Number5[7][11] = 4'hC;
    Number5[8][11] = 4'hC;
    Number5[9][11] = 4'hC;
    Number5[10][11] = 4'hC;
    Number5[11][11] = 4'hC;
    Number5[12][11] = 4'hC;
    Number5[13][11] = 4'hC;
    Number5[14][11] = 4'hD;
    Number5[15][11] = 4'hD;
    Number5[16][11] = 4'hF;
    Number5[17][11] = 4'hF;
    Number5[18][11] = 4'hF;
    Number5[19][11] = 4'hF;
    Number5[20][11] = 4'hF;
    Number5[21][11] = 4'hF;
    Number5[22][11] = 4'hF;
    Number5[0][12] = 4'hF;
    Number5[1][12] = 4'hF;
    Number5[2][12] = 4'hF;
    Number5[3][12] = 4'hF;
    Number5[4][12] = 4'hD;
    Number5[5][12] = 4'hC;
    Number5[6][12] = 4'hC;
    Number5[7][12] = 4'hC;
    Number5[8][12] = 4'hC;
    Number5[9][12] = 4'hC;
    Number5[10][12] = 4'hC;
    Number5[11][12] = 4'hC;
    Number5[12][12] = 4'hC;
    Number5[13][12] = 4'hC;
    Number5[14][12] = 4'hC;
    Number5[15][12] = 4'hC;
    Number5[16][12] = 4'hC;
    Number5[17][12] = 4'hD;
    Number5[18][12] = 4'hF;
    Number5[19][12] = 4'hF;
    Number5[20][12] = 4'hF;
    Number5[21][12] = 4'hF;
    Number5[22][12] = 4'hF;
    Number5[0][13] = 4'hF;
    Number5[1][13] = 4'hF;
    Number5[2][13] = 4'hF;
    Number5[3][13] = 4'hF;
    Number5[4][13] = 4'hD;
    Number5[5][13] = 4'hC;
    Number5[6][13] = 4'hC;
    Number5[7][13] = 4'hC;
    Number5[8][13] = 4'hC;
    Number5[9][13] = 4'hC;
    Number5[10][13] = 4'hC;
    Number5[11][13] = 4'hC;
    Number5[12][13] = 4'hC;
    Number5[13][13] = 4'hC;
    Number5[14][13] = 4'hC;
    Number5[15][13] = 4'hC;
    Number5[16][13] = 4'hC;
    Number5[17][13] = 4'hC;
    Number5[18][13] = 4'hD;
    Number5[19][13] = 4'hF;
    Number5[20][13] = 4'hF;
    Number5[21][13] = 4'hF;
    Number5[22][13] = 4'hF;
    Number5[0][14] = 4'hF;
    Number5[1][14] = 4'hF;
    Number5[2][14] = 4'hF;
    Number5[3][14] = 4'hF;
    Number5[4][14] = 4'hD;
    Number5[5][14] = 4'hC;
    Number5[6][14] = 4'hC;
    Number5[7][14] = 4'hC;
    Number5[8][14] = 4'hC;
    Number5[9][14] = 4'hC;
    Number5[10][14] = 4'hC;
    Number5[11][14] = 4'hC;
    Number5[12][14] = 4'hC;
    Number5[13][14] = 4'hC;
    Number5[14][14] = 4'hC;
    Number5[15][14] = 4'hC;
    Number5[16][14] = 4'hC;
    Number5[17][14] = 4'hC;
    Number5[18][14] = 4'hC;
    Number5[19][14] = 4'hE;
    Number5[20][14] = 4'hF;
    Number5[21][14] = 4'hF;
    Number5[22][14] = 4'hF;
    Number5[0][15] = 4'hF;
    Number5[1][15] = 4'hF;
    Number5[2][15] = 4'hF;
    Number5[3][15] = 4'hF;
    Number5[4][15] = 4'hF;
    Number5[5][15] = 4'hE;
    Number5[6][15] = 4'hE;
    Number5[7][15] = 4'hE;
    Number5[8][15] = 4'hF;
    Number5[9][15] = 4'hF;
    Number5[10][15] = 4'hE;
    Number5[11][15] = 4'hE;
    Number5[12][15] = 4'hD;
    Number5[13][15] = 4'hC;
    Number5[14][15] = 4'hC;
    Number5[15][15] = 4'hC;
    Number5[16][15] = 4'hC;
    Number5[17][15] = 4'hC;
    Number5[18][15] = 4'hC;
    Number5[19][15] = 4'hD;
    Number5[20][15] = 4'hF;
    Number5[21][15] = 4'hF;
    Number5[22][15] = 4'hF;
    Number5[0][16] = 4'hF;
    Number5[1][16] = 4'hF;
    Number5[2][16] = 4'hF;
    Number5[3][16] = 4'hF;
    Number5[4][16] = 4'hF;
    Number5[5][16] = 4'hF;
    Number5[6][16] = 4'hF;
    Number5[7][16] = 4'hF;
    Number5[8][16] = 4'hF;
    Number5[9][16] = 4'hF;
    Number5[10][16] = 4'hF;
    Number5[11][16] = 4'hF;
    Number5[12][16] = 4'hF;
    Number5[13][16] = 4'hD;
    Number5[14][16] = 4'hC;
    Number5[15][16] = 4'hC;
    Number5[16][16] = 4'hC;
    Number5[17][16] = 4'hC;
    Number5[18][16] = 4'hC;
    Number5[19][16] = 4'hC;
    Number5[20][16] = 4'hF;
    Number5[21][16] = 4'hF;
    Number5[22][16] = 4'hF;
    Number5[0][17] = 4'hF;
    Number5[1][17] = 4'hF;
    Number5[2][17] = 4'hF;
    Number5[3][17] = 4'hF;
    Number5[4][17] = 4'hF;
    Number5[5][17] = 4'hF;
    Number5[6][17] = 4'hF;
    Number5[7][17] = 4'hF;
    Number5[8][17] = 4'hF;
    Number5[9][17] = 4'hF;
    Number5[10][17] = 4'hF;
    Number5[11][17] = 4'hF;
    Number5[12][17] = 4'hF;
    Number5[13][17] = 4'hF;
    Number5[14][17] = 4'hC;
    Number5[15][17] = 4'hC;
    Number5[16][17] = 4'hC;
    Number5[17][17] = 4'hC;
    Number5[18][17] = 4'hC;
    Number5[19][17] = 4'hC;
    Number5[20][17] = 4'hF;
    Number5[21][17] = 4'hF;
    Number5[22][17] = 4'hF;
    Number5[0][18] = 4'hF;
    Number5[1][18] = 4'hF;
    Number5[2][18] = 4'hF;
    Number5[3][18] = 4'hF;
    Number5[4][18] = 4'hF;
    Number5[5][18] = 4'hF;
    Number5[6][18] = 4'hF;
    Number5[7][18] = 4'hF;
    Number5[8][18] = 4'hF;
    Number5[9][18] = 4'hF;
    Number5[10][18] = 4'hF;
    Number5[11][18] = 4'hF;
    Number5[12][18] = 4'hF;
    Number5[13][18] = 4'hF;
    Number5[14][18] = 4'hD;
    Number5[15][18] = 4'hC;
    Number5[16][18] = 4'hC;
    Number5[17][18] = 4'hC;
    Number5[18][18] = 4'hC;
    Number5[19][18] = 4'hC;
    Number5[20][18] = 4'hF;
    Number5[21][18] = 4'hF;
    Number5[22][18] = 4'hF;
    Number5[0][19] = 4'hF;
    Number5[1][19] = 4'hF;
    Number5[2][19] = 4'hF;
    Number5[3][19] = 4'hF;
    Number5[4][19] = 4'hF;
    Number5[5][19] = 4'hF;
    Number5[6][19] = 4'hF;
    Number5[7][19] = 4'hF;
    Number5[8][19] = 4'hF;
    Number5[9][19] = 4'hF;
    Number5[10][19] = 4'hF;
    Number5[11][19] = 4'hF;
    Number5[12][19] = 4'hF;
    Number5[13][19] = 4'hF;
    Number5[14][19] = 4'hD;
    Number5[15][19] = 4'hC;
    Number5[16][19] = 4'hC;
    Number5[17][19] = 4'hC;
    Number5[18][19] = 4'hC;
    Number5[19][19] = 4'hC;
    Number5[20][19] = 4'hF;
    Number5[21][19] = 4'hF;
    Number5[22][19] = 4'hF;
    Number5[0][20] = 4'hF;
    Number5[1][20] = 4'hF;
    Number5[2][20] = 4'hF;
    Number5[3][20] = 4'hF;
    Number5[4][20] = 4'hF;
    Number5[5][20] = 4'hF;
    Number5[6][20] = 4'hF;
    Number5[7][20] = 4'hF;
    Number5[8][20] = 4'hF;
    Number5[9][20] = 4'hF;
    Number5[10][20] = 4'hF;
    Number5[11][20] = 4'hF;
    Number5[12][20] = 4'hF;
    Number5[13][20] = 4'hF;
    Number5[14][20] = 4'hC;
    Number5[15][20] = 4'hC;
    Number5[16][20] = 4'hC;
    Number5[17][20] = 4'hC;
    Number5[18][20] = 4'hC;
    Number5[19][20] = 4'hD;
    Number5[20][20] = 4'hF;
    Number5[21][20] = 4'hF;
    Number5[22][20] = 4'hF;
    Number5[0][21] = 4'hF;
    Number5[1][21] = 4'hF;
    Number5[2][21] = 4'hF;
    Number5[3][21] = 4'hF;
    Number5[4][21] = 4'hF;
    Number5[5][21] = 4'hF;
    Number5[6][21] = 4'hF;
    Number5[7][21] = 4'hF;
    Number5[8][21] = 4'hF;
    Number5[9][21] = 4'hF;
    Number5[10][21] = 4'hF;
    Number5[11][21] = 4'hF;
    Number5[12][21] = 4'hF;
    Number5[13][21] = 4'hD;
    Number5[14][21] = 4'hC;
    Number5[15][21] = 4'hC;
    Number5[16][21] = 4'hC;
    Number5[17][21] = 4'hC;
    Number5[18][21] = 4'hC;
    Number5[19][21] = 4'hD;
    Number5[20][21] = 4'hF;
    Number5[21][21] = 4'hF;
    Number5[22][21] = 4'hF;
    Number5[0][22] = 4'hF;
    Number5[1][22] = 4'hF;
    Number5[2][22] = 4'hF;
    Number5[3][22] = 4'hD;
    Number5[4][22] = 4'hC;
    Number5[5][22] = 4'hD;
    Number5[6][22] = 4'hD;
    Number5[7][22] = 4'hE;
    Number5[8][22] = 4'hF;
    Number5[9][22] = 4'hF;
    Number5[10][22] = 4'hE;
    Number5[11][22] = 4'hE;
    Number5[12][22] = 4'hD;
    Number5[13][22] = 4'hC;
    Number5[14][22] = 4'hC;
    Number5[15][22] = 4'hC;
    Number5[16][22] = 4'hC;
    Number5[17][22] = 4'hC;
    Number5[18][22] = 4'hC;
    Number5[19][22] = 4'hF;
    Number5[20][22] = 4'hF;
    Number5[21][22] = 4'hF;
    Number5[22][22] = 4'hF;
    Number5[0][23] = 4'hF;
    Number5[1][23] = 4'hF;
    Number5[2][23] = 4'hF;
    Number5[3][23] = 4'hD;
    Number5[4][23] = 4'hC;
    Number5[5][23] = 4'hC;
    Number5[6][23] = 4'hC;
    Number5[7][23] = 4'hC;
    Number5[8][23] = 4'hC;
    Number5[9][23] = 4'hC;
    Number5[10][23] = 4'hC;
    Number5[11][23] = 4'hC;
    Number5[12][23] = 4'hC;
    Number5[13][23] = 4'hC;
    Number5[14][23] = 4'hC;
    Number5[15][23] = 4'hC;
    Number5[16][23] = 4'hC;
    Number5[17][23] = 4'hC;
    Number5[18][23] = 4'hD;
    Number5[19][23] = 4'hF;
    Number5[20][23] = 4'hF;
    Number5[21][23] = 4'hF;
    Number5[22][23] = 4'hF;
    Number5[0][24] = 4'hF;
    Number5[1][24] = 4'hF;
    Number5[2][24] = 4'hF;
    Number5[3][24] = 4'hD;
    Number5[4][24] = 4'hC;
    Number5[5][24] = 4'hC;
    Number5[6][24] = 4'hC;
    Number5[7][24] = 4'hC;
    Number5[8][24] = 4'hC;
    Number5[9][24] = 4'hC;
    Number5[10][24] = 4'hC;
    Number5[11][24] = 4'hC;
    Number5[12][24] = 4'hC;
    Number5[13][24] = 4'hC;
    Number5[14][24] = 4'hC;
    Number5[15][24] = 4'hC;
    Number5[16][24] = 4'hC;
    Number5[17][24] = 4'hD;
    Number5[18][24] = 4'hF;
    Number5[19][24] = 4'hF;
    Number5[20][24] = 4'hF;
    Number5[21][24] = 4'hF;
    Number5[22][24] = 4'hF;
    Number5[0][25] = 4'hF;
    Number5[1][25] = 4'hF;
    Number5[2][25] = 4'hF;
    Number5[3][25] = 4'hD;
    Number5[4][25] = 4'hC;
    Number5[5][25] = 4'hC;
    Number5[6][25] = 4'hC;
    Number5[7][25] = 4'hC;
    Number5[8][25] = 4'hC;
    Number5[9][25] = 4'hC;
    Number5[10][25] = 4'hC;
    Number5[11][25] = 4'hC;
    Number5[12][25] = 4'hC;
    Number5[13][25] = 4'hC;
    Number5[14][25] = 4'hC;
    Number5[15][25] = 4'hC;
    Number5[16][25] = 4'hE;
    Number5[17][25] = 4'hF;
    Number5[18][25] = 4'hF;
    Number5[19][25] = 4'hF;
    Number5[20][25] = 4'hF;
    Number5[21][25] = 4'hF;
    Number5[22][25] = 4'hF;
    Number5[0][26] = 4'hF;
    Number5[1][26] = 4'hF;
    Number5[2][26] = 4'hF;
    Number5[3][26] = 4'hF;
    Number5[4][26] = 4'hE;
    Number5[5][26] = 4'hD;
    Number5[6][26] = 4'hD;
    Number5[7][26] = 4'hC;
    Number5[8][26] = 4'hC;
    Number5[9][26] = 4'hC;
    Number5[10][26] = 4'hC;
    Number5[11][26] = 4'hC;
    Number5[12][26] = 4'hC;
    Number5[13][26] = 4'hD;
    Number5[14][26] = 4'hE;
    Number5[15][26] = 4'hF;
    Number5[16][26] = 4'hF;
    Number5[17][26] = 4'hF;
    Number5[18][26] = 4'hF;
    Number5[19][26] = 4'hF;
    Number5[20][26] = 4'hF;
    Number5[21][26] = 4'hF;
    Number5[22][26] = 4'hF;
    Number5[0][27] = 4'hF;
    Number5[1][27] = 4'hF;
    Number5[2][27] = 4'hF;
    Number5[3][27] = 4'hF;
    Number5[4][27] = 4'hF;
    Number5[5][27] = 4'hF;
    Number5[6][27] = 4'hF;
    Number5[7][27] = 4'hF;
    Number5[8][27] = 4'hF;
    Number5[9][27] = 4'hF;
    Number5[10][27] = 4'hF;
    Number5[11][27] = 4'hF;
    Number5[12][27] = 4'hF;
    Number5[13][27] = 4'hF;
    Number5[14][27] = 4'hF;
    Number5[15][27] = 4'hF;
    Number5[16][27] = 4'hF;
    Number5[17][27] = 4'hF;
    Number5[18][27] = 4'hF;
    Number5[19][27] = 4'hF;
    Number5[20][27] = 4'hF;
    Number5[21][27] = 4'hF;
    Number5[22][27] = 4'hF;
    Number5[0][28] = 4'hF;
    Number5[1][28] = 4'hF;
    Number5[2][28] = 4'hF;
    Number5[3][28] = 4'hF;
    Number5[4][28] = 4'hF;
    Number5[5][28] = 4'hF;
    Number5[6][28] = 4'hF;
    Number5[7][28] = 4'hF;
    Number5[8][28] = 4'hF;
    Number5[9][28] = 4'hF;
    Number5[10][28] = 4'hF;
    Number5[11][28] = 4'hF;
    Number5[12][28] = 4'hF;
    Number5[13][28] = 4'hF;
    Number5[14][28] = 4'hF;
    Number5[15][28] = 4'hF;
    Number5[16][28] = 4'hF;
    Number5[17][28] = 4'hF;
    Number5[18][28] = 4'hF;
    Number5[19][28] = 4'hF;
    Number5[20][28] = 4'hF;
    Number5[21][28] = 4'hF;
    Number5[22][28] = 4'hF;

// Number 6
    Number6[0][0] = 4'hF;
    Number6[1][0] = 4'hF;
    Number6[2][0] = 4'hF;
    Number6[3][0] = 4'hF;
    Number6[4][0] = 4'hF;
    Number6[5][0] = 4'hF;
    Number6[6][0] = 4'hF;
    Number6[7][0] = 4'hF;
    Number6[8][0] = 4'hF;
    Number6[9][0] = 4'hF;
    Number6[10][0] = 4'hF;
    Number6[11][0] = 4'hF;
    Number6[12][0] = 4'hF;
    Number6[13][0] = 4'hF;
    Number6[14][0] = 4'hF;
    Number6[15][0] = 4'hF;
    Number6[16][0] = 4'hF;
    Number6[17][0] = 4'hF;
    Number6[18][0] = 4'hF;
    Number6[19][0] = 4'hF;
    Number6[20][0] = 4'hF;
    Number6[21][0] = 4'hF;
    Number6[22][0] = 4'hF;
    Number6[0][1] = 4'hF;
    Number6[1][1] = 4'hF;
    Number6[2][1] = 4'hF;
    Number6[3][1] = 4'hF;
    Number6[4][1] = 4'hF;
    Number6[5][1] = 4'hF;
    Number6[6][1] = 4'hF;
    Number6[7][1] = 4'hF;
    Number6[8][1] = 4'hF;
    Number6[9][1] = 4'hF;
    Number6[10][1] = 4'hF;
    Number6[11][1] = 4'hF;
    Number6[12][1] = 4'hF;
    Number6[13][1] = 4'hF;
    Number6[14][1] = 4'hF;
    Number6[15][1] = 4'hF;
    Number6[16][1] = 4'hF;
    Number6[17][1] = 4'hF;
    Number6[18][1] = 4'hF;
    Number6[19][1] = 4'hF;
    Number6[20][1] = 4'hF;
    Number6[21][1] = 4'hF;
    Number6[22][1] = 4'hF;
    Number6[0][2] = 4'hF;
    Number6[1][2] = 4'hF;
    Number6[2][2] = 4'hF;
    Number6[3][2] = 4'hF;
    Number6[4][2] = 4'hF;
    Number6[5][2] = 4'hF;
    Number6[6][2] = 4'hF;
    Number6[7][2] = 4'hF;
    Number6[8][2] = 4'hF;
    Number6[9][2] = 4'hE;
    Number6[10][2] = 4'hD;
    Number6[11][2] = 4'hC;
    Number6[12][2] = 4'hC;
    Number6[13][2] = 4'hC;
    Number6[14][2] = 4'hC;
    Number6[15][2] = 4'hC;
    Number6[16][2] = 4'hC;
    Number6[17][2] = 4'hD;
    Number6[18][2] = 4'hE;
    Number6[19][2] = 4'hF;
    Number6[20][2] = 4'hF;
    Number6[21][2] = 4'hF;
    Number6[22][2] = 4'hF;
    Number6[0][3] = 4'hF;
    Number6[1][3] = 4'hF;
    Number6[2][3] = 4'hF;
    Number6[3][3] = 4'hF;
    Number6[4][3] = 4'hF;
    Number6[5][3] = 4'hF;
    Number6[6][3] = 4'hF;
    Number6[7][3] = 4'hE;
    Number6[8][3] = 4'hC;
    Number6[9][3] = 4'hC;
    Number6[10][3] = 4'hC;
    Number6[11][3] = 4'hC;
    Number6[12][3] = 4'hC;
    Number6[13][3] = 4'hC;
    Number6[14][3] = 4'hC;
    Number6[15][3] = 4'hC;
    Number6[16][3] = 4'hC;
    Number6[17][3] = 4'hC;
    Number6[18][3] = 4'hC;
    Number6[19][3] = 4'hF;
    Number6[20][3] = 4'hF;
    Number6[21][3] = 4'hF;
    Number6[22][3] = 4'hF;
    Number6[0][4] = 4'hF;
    Number6[1][4] = 4'hF;
    Number6[2][4] = 4'hF;
    Number6[3][4] = 4'hF;
    Number6[4][4] = 4'hF;
    Number6[5][4] = 4'hF;
    Number6[6][4] = 4'hD;
    Number6[7][4] = 4'hC;
    Number6[8][4] = 4'hC;
    Number6[9][4] = 4'hC;
    Number6[10][4] = 4'hC;
    Number6[11][4] = 4'hC;
    Number6[12][4] = 4'hC;
    Number6[13][4] = 4'hC;
    Number6[14][4] = 4'hC;
    Number6[15][4] = 4'hC;
    Number6[16][4] = 4'hC;
    Number6[17][4] = 4'hC;
    Number6[18][4] = 4'hC;
    Number6[19][4] = 4'hF;
    Number6[20][4] = 4'hF;
    Number6[21][4] = 4'hF;
    Number6[22][4] = 4'hF;
    Number6[0][5] = 4'hF;
    Number6[1][5] = 4'hF;
    Number6[2][5] = 4'hF;
    Number6[3][5] = 4'hF;
    Number6[4][5] = 4'hF;
    Number6[5][5] = 4'hE;
    Number6[6][5] = 4'hC;
    Number6[7][5] = 4'hC;
    Number6[8][5] = 4'hC;
    Number6[9][5] = 4'hC;
    Number6[10][5] = 4'hC;
    Number6[11][5] = 4'hC;
    Number6[12][5] = 4'hC;
    Number6[13][5] = 4'hC;
    Number6[14][5] = 4'hC;
    Number6[15][5] = 4'hC;
    Number6[16][5] = 4'hC;
    Number6[17][5] = 4'hC;
    Number6[18][5] = 4'hC;
    Number6[19][5] = 4'hF;
    Number6[20][5] = 4'hF;
    Number6[21][5] = 4'hF;
    Number6[22][5] = 4'hF;
    Number6[0][6] = 4'hF;
    Number6[1][6] = 4'hF;
    Number6[2][6] = 4'hF;
    Number6[3][6] = 4'hF;
    Number6[4][6] = 4'hF;
    Number6[5][6] = 4'hC;
    Number6[6][6] = 4'hC;
    Number6[7][6] = 4'hC;
    Number6[8][6] = 4'hC;
    Number6[9][6] = 4'hC;
    Number6[10][6] = 4'hC;
    Number6[11][6] = 4'hD;
    Number6[12][6] = 4'hE;
    Number6[13][6] = 4'hF;
    Number6[14][6] = 4'hF;
    Number6[15][6] = 4'hE;
    Number6[16][6] = 4'hD;
    Number6[17][6] = 4'hD;
    Number6[18][6] = 4'hD;
    Number6[19][6] = 4'hF;
    Number6[20][6] = 4'hF;
    Number6[21][6] = 4'hF;
    Number6[22][6] = 4'hF;
    Number6[0][7] = 4'hF;
    Number6[1][7] = 4'hF;
    Number6[2][7] = 4'hF;
    Number6[3][7] = 4'hF;
    Number6[4][7] = 4'hD;
    Number6[5][7] = 4'hC;
    Number6[6][7] = 4'hC;
    Number6[7][7] = 4'hC;
    Number6[8][7] = 4'hC;
    Number6[9][7] = 4'hC;
    Number6[10][7] = 4'hE;
    Number6[11][7] = 4'hF;
    Number6[12][7] = 4'hF;
    Number6[13][7] = 4'hF;
    Number6[14][7] = 4'hF;
    Number6[15][7] = 4'hF;
    Number6[16][7] = 4'hF;
    Number6[17][7] = 4'hF;
    Number6[18][7] = 4'hF;
    Number6[19][7] = 4'hF;
    Number6[20][7] = 4'hF;
    Number6[21][7] = 4'hF;
    Number6[22][7] = 4'hF;
    Number6[0][8] = 4'hF;
    Number6[1][8] = 4'hF;
    Number6[2][8] = 4'hF;
    Number6[3][8] = 4'hF;
    Number6[4][8] = 4'hC;
    Number6[5][8] = 4'hC;
    Number6[6][8] = 4'hC;
    Number6[7][8] = 4'hC;
    Number6[8][8] = 4'hC;
    Number6[9][8] = 4'hE;
    Number6[10][8] = 4'hF;
    Number6[11][8] = 4'hF;
    Number6[12][8] = 4'hF;
    Number6[13][8] = 4'hF;
    Number6[14][8] = 4'hF;
    Number6[15][8] = 4'hF;
    Number6[16][8] = 4'hF;
    Number6[17][8] = 4'hF;
    Number6[18][8] = 4'hF;
    Number6[19][8] = 4'hF;
    Number6[20][8] = 4'hF;
    Number6[21][8] = 4'hF;
    Number6[22][8] = 4'hF;
    Number6[0][9] = 4'hF;
    Number6[1][9] = 4'hF;
    Number6[2][9] = 4'hF;
    Number6[3][9] = 4'hE;
    Number6[4][9] = 4'hC;
    Number6[5][9] = 4'hC;
    Number6[6][9] = 4'hC;
    Number6[7][9] = 4'hC;
    Number6[8][9] = 4'hD;
    Number6[9][9] = 4'hF;
    Number6[10][9] = 4'hF;
    Number6[11][9] = 4'hF;
    Number6[12][9] = 4'hF;
    Number6[13][9] = 4'hF;
    Number6[14][9] = 4'hF;
    Number6[15][9] = 4'hF;
    Number6[16][9] = 4'hF;
    Number6[17][9] = 4'hF;
    Number6[18][9] = 4'hF;
    Number6[19][9] = 4'hF;
    Number6[20][9] = 4'hF;
    Number6[21][9] = 4'hF;
    Number6[22][9] = 4'hF;
    Number6[0][10] = 4'hF;
    Number6[1][10] = 4'hF;
    Number6[2][10] = 4'hF;
    Number6[3][10] = 4'hD;
    Number6[4][10] = 4'hC;
    Number6[5][10] = 4'hC;
    Number6[6][10] = 4'hC;
    Number6[7][10] = 4'hC;
    Number6[8][10] = 4'hD;
    Number6[9][10] = 4'hF;
    Number6[10][10] = 4'hF;
    Number6[11][10] = 4'hF;
    Number6[12][10] = 4'hF;
    Number6[13][10] = 4'hF;
    Number6[14][10] = 4'hF;
    Number6[15][10] = 4'hF;
    Number6[16][10] = 4'hF;
    Number6[17][10] = 4'hF;
    Number6[18][10] = 4'hF;
    Number6[19][10] = 4'hF;
    Number6[20][10] = 4'hF;
    Number6[21][10] = 4'hF;
    Number6[22][10] = 4'hF;
    Number6[0][11] = 4'hF;
    Number6[1][11] = 4'hF;
    Number6[2][11] = 4'hF;
    Number6[3][11] = 4'hD;
    Number6[4][11] = 4'hC;
    Number6[5][11] = 4'hC;
    Number6[6][11] = 4'hC;
    Number6[7][11] = 4'hC;
    Number6[8][11] = 4'hE;
    Number6[9][11] = 4'hE;
    Number6[10][11] = 4'hD;
    Number6[11][11] = 4'hC;
    Number6[12][11] = 4'hC;
    Number6[13][11] = 4'hC;
    Number6[14][11] = 4'hC;
    Number6[15][11] = 4'hC;
    Number6[16][11] = 4'hD;
    Number6[17][11] = 4'hE;
    Number6[18][11] = 4'hF;
    Number6[19][11] = 4'hF;
    Number6[20][11] = 4'hF;
    Number6[21][11] = 4'hF;
    Number6[22][11] = 4'hF;
    Number6[0][12] = 4'hF;
    Number6[1][12] = 4'hF;
    Number6[2][12] = 4'hF;
    Number6[3][12] = 4'hC;
    Number6[4][12] = 4'hC;
    Number6[5][12] = 4'hC;
    Number6[6][12] = 4'hC;
    Number6[7][12] = 4'hC;
    Number6[8][12] = 4'hC;
    Number6[9][12] = 4'hC;
    Number6[10][12] = 4'hC;
    Number6[11][12] = 4'hC;
    Number6[12][12] = 4'hC;
    Number6[13][12] = 4'hC;
    Number6[14][12] = 4'hC;
    Number6[15][12] = 4'hC;
    Number6[16][12] = 4'hC;
    Number6[17][12] = 4'hC;
    Number6[18][12] = 4'hD;
    Number6[19][12] = 4'hF;
    Number6[20][12] = 4'hF;
    Number6[21][12] = 4'hF;
    Number6[22][12] = 4'hF;
    Number6[0][13] = 4'hF;
    Number6[1][13] = 4'hF;
    Number6[2][13] = 4'hF;
    Number6[3][13] = 4'hC;
    Number6[4][13] = 4'hC;
    Number6[5][13] = 4'hC;
    Number6[6][13] = 4'hC;
    Number6[7][13] = 4'hC;
    Number6[8][13] = 4'hC;
    Number6[9][13] = 4'hC;
    Number6[10][13] = 4'hC;
    Number6[11][13] = 4'hC;
    Number6[12][13] = 4'hC;
    Number6[13][13] = 4'hC;
    Number6[14][13] = 4'hC;
    Number6[15][13] = 4'hC;
    Number6[16][13] = 4'hC;
    Number6[17][13] = 4'hC;
    Number6[18][13] = 4'hC;
    Number6[19][13] = 4'hD;
    Number6[20][13] = 4'hF;
    Number6[21][13] = 4'hF;
    Number6[22][13] = 4'hF;
    Number6[0][14] = 4'hF;
    Number6[1][14] = 4'hF;
    Number6[2][14] = 4'hF;
    Number6[3][14] = 4'hC;
    Number6[4][14] = 4'hC;
    Number6[5][14] = 4'hC;
    Number6[6][14] = 4'hC;
    Number6[7][14] = 4'hC;
    Number6[8][14] = 4'hC;
    Number6[9][14] = 4'hC;
    Number6[10][14] = 4'hC;
    Number6[11][14] = 4'hC;
    Number6[12][14] = 4'hC;
    Number6[13][14] = 4'hC;
    Number6[14][14] = 4'hC;
    Number6[15][14] = 4'hC;
    Number6[16][14] = 4'hC;
    Number6[17][14] = 4'hC;
    Number6[18][14] = 4'hC;
    Number6[19][14] = 4'hC;
    Number6[20][14] = 4'hF;
    Number6[21][14] = 4'hF;
    Number6[22][14] = 4'hF;
    Number6[0][15] = 4'hF;
    Number6[1][15] = 4'hF;
    Number6[2][15] = 4'hF;
    Number6[3][15] = 4'hC;
    Number6[4][15] = 4'hC;
    Number6[5][15] = 4'hC;
    Number6[6][15] = 4'hC;
    Number6[7][15] = 4'hC;
    Number6[8][15] = 4'hC;
    Number6[9][15] = 4'hD;
    Number6[10][15] = 4'hD;
    Number6[11][15] = 4'hE;
    Number6[12][15] = 4'hF;
    Number6[13][15] = 4'hE;
    Number6[14][15] = 4'hC;
    Number6[15][15] = 4'hC;
    Number6[16][15] = 4'hC;
    Number6[17][15] = 4'hC;
    Number6[18][15] = 4'hC;
    Number6[19][15] = 4'hC;
    Number6[20][15] = 4'hE;
    Number6[21][15] = 4'hF;
    Number6[22][15] = 4'hF;
    Number6[0][16] = 4'hF;
    Number6[1][16] = 4'hF;
    Number6[2][16] = 4'hF;
    Number6[3][16] = 4'hC;
    Number6[4][16] = 4'hC;
    Number6[5][16] = 4'hC;
    Number6[6][16] = 4'hC;
    Number6[7][16] = 4'hC;
    Number6[8][16] = 4'hD;
    Number6[9][16] = 4'hF;
    Number6[10][16] = 4'hF;
    Number6[11][16] = 4'hF;
    Number6[12][16] = 4'hF;
    Number6[13][16] = 4'hF;
    Number6[14][16] = 4'hF;
    Number6[15][16] = 4'hC;
    Number6[16][16] = 4'hC;
    Number6[17][16] = 4'hC;
    Number6[18][16] = 4'hC;
    Number6[19][16] = 4'hC;
    Number6[20][16] = 4'hD;
    Number6[21][16] = 4'hF;
    Number6[22][16] = 4'hF;
    Number6[0][17] = 4'hF;
    Number6[1][17] = 4'hF;
    Number6[2][17] = 4'hF;
    Number6[3][17] = 4'hC;
    Number6[4][17] = 4'hC;
    Number6[5][17] = 4'hC;
    Number6[6][17] = 4'hC;
    Number6[7][17] = 4'hC;
    Number6[8][17] = 4'hD;
    Number6[9][17] = 4'hF;
    Number6[10][17] = 4'hF;
    Number6[11][17] = 4'hF;
    Number6[12][17] = 4'hF;
    Number6[13][17] = 4'hF;
    Number6[14][17] = 4'hF;
    Number6[15][17] = 4'hD;
    Number6[16][17] = 4'hC;
    Number6[17][17] = 4'hC;
    Number6[18][17] = 4'hC;
    Number6[19][17] = 4'hC;
    Number6[20][17] = 4'hD;
    Number6[21][17] = 4'hF;
    Number6[22][17] = 4'hF;
    Number6[0][18] = 4'hF;
    Number6[1][18] = 4'hF;
    Number6[2][18] = 4'hF;
    Number6[3][18] = 4'hC;
    Number6[4][18] = 4'hC;
    Number6[5][18] = 4'hC;
    Number6[6][18] = 4'hC;
    Number6[7][18] = 4'hC;
    Number6[8][18] = 4'hD;
    Number6[9][18] = 4'hF;
    Number6[10][18] = 4'hF;
    Number6[11][18] = 4'hF;
    Number6[12][18] = 4'hF;
    Number6[13][18] = 4'hF;
    Number6[14][18] = 4'hF;
    Number6[15][18] = 4'hD;
    Number6[16][18] = 4'hC;
    Number6[17][18] = 4'hC;
    Number6[18][18] = 4'hC;
    Number6[19][18] = 4'hC;
    Number6[20][18] = 4'hD;
    Number6[21][18] = 4'hF;
    Number6[22][18] = 4'hF;
    Number6[0][19] = 4'hF;
    Number6[1][19] = 4'hF;
    Number6[2][19] = 4'hF;
    Number6[3][19] = 4'hD;
    Number6[4][19] = 4'hC;
    Number6[5][19] = 4'hC;
    Number6[6][19] = 4'hC;
    Number6[7][19] = 4'hC;
    Number6[8][19] = 4'hD;
    Number6[9][19] = 4'hF;
    Number6[10][19] = 4'hF;
    Number6[11][19] = 4'hF;
    Number6[12][19] = 4'hF;
    Number6[13][19] = 4'hF;
    Number6[14][19] = 4'hF;
    Number6[15][19] = 4'hD;
    Number6[16][19] = 4'hC;
    Number6[17][19] = 4'hC;
    Number6[18][19] = 4'hC;
    Number6[19][19] = 4'hC;
    Number6[20][19] = 4'hD;
    Number6[21][19] = 4'hF;
    Number6[22][19] = 4'hF;
    Number6[0][20] = 4'hF;
    Number6[1][20] = 4'hF;
    Number6[2][20] = 4'hF;
    Number6[3][20] = 4'hD;
    Number6[4][20] = 4'hC;
    Number6[5][20] = 4'hC;
    Number6[6][20] = 4'hC;
    Number6[7][20] = 4'hC;
    Number6[8][20] = 4'hC;
    Number6[9][20] = 4'hF;
    Number6[10][20] = 4'hF;
    Number6[11][20] = 4'hF;
    Number6[12][20] = 4'hF;
    Number6[13][20] = 4'hF;
    Number6[14][20] = 4'hF;
    Number6[15][20] = 4'hC;
    Number6[16][20] = 4'hC;
    Number6[17][20] = 4'hC;
    Number6[18][20] = 4'hC;
    Number6[19][20] = 4'hC;
    Number6[20][20] = 4'hD;
    Number6[21][20] = 4'hF;
    Number6[22][20] = 4'hF;
    Number6[0][21] = 4'hF;
    Number6[1][21] = 4'hF;
    Number6[2][21] = 4'hF;
    Number6[3][21] = 4'hE;
    Number6[4][21] = 4'hC;
    Number6[5][21] = 4'hC;
    Number6[6][21] = 4'hC;
    Number6[7][21] = 4'hC;
    Number6[8][21] = 4'hC;
    Number6[9][21] = 4'hE;
    Number6[10][21] = 4'hF;
    Number6[11][21] = 4'hF;
    Number6[12][21] = 4'hF;
    Number6[13][21] = 4'hF;
    Number6[14][21] = 4'hE;
    Number6[15][21] = 4'hC;
    Number6[16][21] = 4'hC;
    Number6[17][21] = 4'hC;
    Number6[18][21] = 4'hC;
    Number6[19][21] = 4'hC;
    Number6[20][21] = 4'hE;
    Number6[21][21] = 4'hF;
    Number6[22][21] = 4'hF;
    Number6[0][22] = 4'hF;
    Number6[1][22] = 4'hF;
    Number6[2][22] = 4'hF;
    Number6[3][22] = 4'hF;
    Number6[4][22] = 4'hC;
    Number6[5][22] = 4'hC;
    Number6[6][22] = 4'hC;
    Number6[7][22] = 4'hC;
    Number6[8][22] = 4'hC;
    Number6[9][22] = 4'hC;
    Number6[10][22] = 4'hD;
    Number6[11][22] = 4'hF;
    Number6[12][22] = 4'hE;
    Number6[13][22] = 4'hD;
    Number6[14][22] = 4'hC;
    Number6[15][22] = 4'hC;
    Number6[16][22] = 4'hC;
    Number6[17][22] = 4'hC;
    Number6[18][22] = 4'hC;
    Number6[19][22] = 4'hD;
    Number6[20][22] = 4'hF;
    Number6[21][22] = 4'hF;
    Number6[22][22] = 4'hF;
    Number6[0][23] = 4'hF;
    Number6[1][23] = 4'hF;
    Number6[2][23] = 4'hF;
    Number6[3][23] = 4'hF;
    Number6[4][23] = 4'hD;
    Number6[5][23] = 4'hC;
    Number6[6][23] = 4'hC;
    Number6[7][23] = 4'hC;
    Number6[8][23] = 4'hC;
    Number6[9][23] = 4'hC;
    Number6[10][23] = 4'hC;
    Number6[11][23] = 4'hC;
    Number6[12][23] = 4'hC;
    Number6[13][23] = 4'hC;
    Number6[14][23] = 4'hC;
    Number6[15][23] = 4'hC;
    Number6[16][23] = 4'hC;
    Number6[17][23] = 4'hC;
    Number6[18][23] = 4'hC;
    Number6[19][23] = 4'hE;
    Number6[20][23] = 4'hF;
    Number6[21][23] = 4'hF;
    Number6[22][23] = 4'hF;
    Number6[0][24] = 4'hF;
    Number6[1][24] = 4'hF;
    Number6[2][24] = 4'hF;
    Number6[3][24] = 4'hF;
    Number6[4][24] = 4'hF;
    Number6[5][24] = 4'hC;
    Number6[6][24] = 4'hC;
    Number6[7][24] = 4'hC;
    Number6[8][24] = 4'hC;
    Number6[9][24] = 4'hC;
    Number6[10][24] = 4'hC;
    Number6[11][24] = 4'hC;
    Number6[12][24] = 4'hC;
    Number6[13][24] = 4'hC;
    Number6[14][24] = 4'hC;
    Number6[15][24] = 4'hC;
    Number6[16][24] = 4'hC;
    Number6[17][24] = 4'hC;
    Number6[18][24] = 4'hD;
    Number6[19][24] = 4'hF;
    Number6[20][24] = 4'hF;
    Number6[21][24] = 4'hF;
    Number6[22][24] = 4'hF;
    Number6[0][25] = 4'hF;
    Number6[1][25] = 4'hF;
    Number6[2][25] = 4'hF;
    Number6[3][25] = 4'hF;
    Number6[4][25] = 4'hF;
    Number6[5][25] = 4'hF;
    Number6[6][25] = 4'hD;
    Number6[7][25] = 4'hC;
    Number6[8][25] = 4'hC;
    Number6[9][25] = 4'hC;
    Number6[10][25] = 4'hC;
    Number6[11][25] = 4'hC;
    Number6[12][25] = 4'hC;
    Number6[13][25] = 4'hC;
    Number6[14][25] = 4'hC;
    Number6[15][25] = 4'hC;
    Number6[16][25] = 4'hC;
    Number6[17][25] = 4'hE;
    Number6[18][25] = 4'hF;
    Number6[19][25] = 4'hF;
    Number6[20][25] = 4'hF;
    Number6[21][25] = 4'hF;
    Number6[22][25] = 4'hF;
    Number6[0][26] = 4'hF;
    Number6[1][26] = 4'hF;
    Number6[2][26] = 4'hF;
    Number6[3][26] = 4'hF;
    Number6[4][26] = 4'hF;
    Number6[5][26] = 4'hF;
    Number6[6][26] = 4'hF;
    Number6[7][26] = 4'hE;
    Number6[8][26] = 4'hD;
    Number6[9][26] = 4'hC;
    Number6[10][26] = 4'hC;
    Number6[11][26] = 4'hC;
    Number6[12][26] = 4'hC;
    Number6[13][26] = 4'hC;
    Number6[14][26] = 4'hD;
    Number6[15][26] = 4'hD;
    Number6[16][26] = 4'hF;
    Number6[17][26] = 4'hF;
    Number6[18][26] = 4'hF;
    Number6[19][26] = 4'hF;
    Number6[20][26] = 4'hF;
    Number6[21][26] = 4'hF;
    Number6[22][26] = 4'hF;
    Number6[0][27] = 4'hF;
    Number6[1][27] = 4'hF;
    Number6[2][27] = 4'hF;
    Number6[3][27] = 4'hF;
    Number6[4][27] = 4'hF;
    Number6[5][27] = 4'hF;
    Number6[6][27] = 4'hF;
    Number6[7][27] = 4'hF;
    Number6[8][27] = 4'hF;
    Number6[9][27] = 4'hF;
    Number6[10][27] = 4'hF;
    Number6[11][27] = 4'hF;
    Number6[12][27] = 4'hF;
    Number6[13][27] = 4'hF;
    Number6[14][27] = 4'hF;
    Number6[15][27] = 4'hF;
    Number6[16][27] = 4'hF;
    Number6[17][27] = 4'hF;
    Number6[18][27] = 4'hF;
    Number6[19][27] = 4'hF;
    Number6[20][27] = 4'hF;
    Number6[21][27] = 4'hF;
    Number6[22][27] = 4'hF;
    Number6[0][28] = 4'hF;
    Number6[1][28] = 4'hF;
    Number6[2][28] = 4'hF;
    Number6[3][28] = 4'hF;
    Number6[4][28] = 4'hF;
    Number6[5][28] = 4'hF;
    Number6[6][28] = 4'hF;
    Number6[7][28] = 4'hF;
    Number6[8][28] = 4'hF;
    Number6[9][28] = 4'hF;
    Number6[10][28] = 4'hF;
    Number6[11][28] = 4'hF;
    Number6[12][28] = 4'hF;
    Number6[13][28] = 4'hF;
    Number6[14][28] = 4'hF;
    Number6[15][28] = 4'hF;
    Number6[16][28] = 4'hF;
    Number6[17][28] = 4'hF;
    Number6[18][28] = 4'hF;
    Number6[19][28] = 4'hF;
    Number6[20][28] = 4'hF;
    Number6[21][28] = 4'hF;
    Number6[22][28] = 4'hF;

// Number 7
    Number7[0][0] = 4'hF;
    Number7[1][0] = 4'hF;
    Number7[2][0] = 4'hF;
    Number7[3][0] = 4'hF;
    Number7[4][0] = 4'hF;
    Number7[5][0] = 4'hF;
    Number7[6][0] = 4'hF;
    Number7[7][0] = 4'hF;
    Number7[8][0] = 4'hF;
    Number7[9][0] = 4'hF;
    Number7[10][0] = 4'hF;
    Number7[11][0] = 4'hF;
    Number7[12][0] = 4'hF;
    Number7[13][0] = 4'hF;
    Number7[14][0] = 4'hF;
    Number7[15][0] = 4'hF;
    Number7[16][0] = 4'hF;
    Number7[17][0] = 4'hF;
    Number7[18][0] = 4'hF;
    Number7[19][0] = 4'hF;
    Number7[20][0] = 4'hF;
    Number7[21][0] = 4'hF;
    Number7[22][0] = 4'hF;
    Number7[0][1] = 4'hF;
    Number7[1][1] = 4'hF;
    Number7[2][1] = 4'hF;
    Number7[3][1] = 4'hF;
    Number7[4][1] = 4'hF;
    Number7[5][1] = 4'hF;
    Number7[6][1] = 4'hF;
    Number7[7][1] = 4'hF;
    Number7[8][1] = 4'hF;
    Number7[9][1] = 4'hF;
    Number7[10][1] = 4'hF;
    Number7[11][1] = 4'hF;
    Number7[12][1] = 4'hF;
    Number7[13][1] = 4'hF;
    Number7[14][1] = 4'hF;
    Number7[15][1] = 4'hF;
    Number7[16][1] = 4'hF;
    Number7[17][1] = 4'hF;
    Number7[18][1] = 4'hF;
    Number7[19][1] = 4'hF;
    Number7[20][1] = 4'hF;
    Number7[21][1] = 4'hF;
    Number7[22][1] = 4'hF;
    Number7[0][2] = 4'hF;
    Number7[1][2] = 4'hF;
    Number7[2][2] = 4'hF;
    Number7[3][2] = 4'hD;
    Number7[4][2] = 4'hC;
    Number7[5][2] = 4'hC;
    Number7[6][2] = 4'hC;
    Number7[7][2] = 4'hC;
    Number7[8][2] = 4'hC;
    Number7[9][2] = 4'hC;
    Number7[10][2] = 4'hC;
    Number7[11][2] = 4'hC;
    Number7[12][2] = 4'hC;
    Number7[13][2] = 4'hC;
    Number7[14][2] = 4'hC;
    Number7[15][2] = 4'hC;
    Number7[16][2] = 4'hC;
    Number7[17][2] = 4'hC;
    Number7[18][2] = 4'hC;
    Number7[19][2] = 4'hC;
    Number7[20][2] = 4'hF;
    Number7[21][2] = 4'hF;
    Number7[22][2] = 4'hF;
    Number7[0][3] = 4'hF;
    Number7[1][3] = 4'hF;
    Number7[2][3] = 4'hF;
    Number7[3][3] = 4'hC;
    Number7[4][3] = 4'hC;
    Number7[5][3] = 4'hC;
    Number7[6][3] = 4'hC;
    Number7[7][3] = 4'hC;
    Number7[8][3] = 4'hC;
    Number7[9][3] = 4'hC;
    Number7[10][3] = 4'hC;
    Number7[11][3] = 4'hC;
    Number7[12][3] = 4'hC;
    Number7[13][3] = 4'hC;
    Number7[14][3] = 4'hC;
    Number7[15][3] = 4'hC;
    Number7[16][3] = 4'hC;
    Number7[17][3] = 4'hC;
    Number7[18][3] = 4'hC;
    Number7[19][3] = 4'hC;
    Number7[20][3] = 4'hE;
    Number7[21][3] = 4'hF;
    Number7[22][3] = 4'hF;
    Number7[0][4] = 4'hF;
    Number7[1][4] = 4'hF;
    Number7[2][4] = 4'hF;
    Number7[3][4] = 4'hC;
    Number7[4][4] = 4'hC;
    Number7[5][4] = 4'hC;
    Number7[6][4] = 4'hC;
    Number7[7][4] = 4'hC;
    Number7[8][4] = 4'hC;
    Number7[9][4] = 4'hC;
    Number7[10][4] = 4'hC;
    Number7[11][4] = 4'hC;
    Number7[12][4] = 4'hC;
    Number7[13][4] = 4'hC;
    Number7[14][4] = 4'hC;
    Number7[15][4] = 4'hC;
    Number7[16][4] = 4'hC;
    Number7[17][4] = 4'hC;
    Number7[18][4] = 4'hC;
    Number7[19][4] = 4'hC;
    Number7[20][4] = 4'hE;
    Number7[21][4] = 4'hF;
    Number7[22][4] = 4'hF;
    Number7[0][5] = 4'hF;
    Number7[1][5] = 4'hF;
    Number7[2][5] = 4'hF;
    Number7[3][5] = 4'hD;
    Number7[4][5] = 4'hC;
    Number7[5][5] = 4'hC;
    Number7[6][5] = 4'hC;
    Number7[7][5] = 4'hC;
    Number7[8][5] = 4'hC;
    Number7[9][5] = 4'hC;
    Number7[10][5] = 4'hC;
    Number7[11][5] = 4'hC;
    Number7[12][5] = 4'hC;
    Number7[13][5] = 4'hC;
    Number7[14][5] = 4'hC;
    Number7[15][5] = 4'hC;
    Number7[16][5] = 4'hC;
    Number7[17][5] = 4'hC;
    Number7[18][5] = 4'hC;
    Number7[19][5] = 4'hC;
    Number7[20][5] = 4'hF;
    Number7[21][5] = 4'hF;
    Number7[22][5] = 4'hF;
    Number7[0][6] = 4'hF;
    Number7[1][6] = 4'hF;
    Number7[2][6] = 4'hF;
    Number7[3][6] = 4'hF;
    Number7[4][6] = 4'hF;
    Number7[5][6] = 4'hF;
    Number7[6][6] = 4'hF;
    Number7[7][6] = 4'hF;
    Number7[8][6] = 4'hF;
    Number7[9][6] = 4'hF;
    Number7[10][6] = 4'hF;
    Number7[11][6] = 4'hF;
    Number7[12][6] = 4'hF;
    Number7[13][6] = 4'hF;
    Number7[14][6] = 4'hC;
    Number7[15][6] = 4'hC;
    Number7[16][6] = 4'hC;
    Number7[17][6] = 4'hC;
    Number7[18][6] = 4'hC;
    Number7[19][6] = 4'hC;
    Number7[20][6] = 4'hF;
    Number7[21][6] = 4'hF;
    Number7[22][6] = 4'hF;
    Number7[0][7] = 4'hF;
    Number7[1][7] = 4'hF;
    Number7[2][7] = 4'hF;
    Number7[3][7] = 4'hF;
    Number7[4][7] = 4'hF;
    Number7[5][7] = 4'hF;
    Number7[6][7] = 4'hF;
    Number7[7][7] = 4'hF;
    Number7[8][7] = 4'hF;
    Number7[9][7] = 4'hF;
    Number7[10][7] = 4'hF;
    Number7[11][7] = 4'hF;
    Number7[12][7] = 4'hF;
    Number7[13][7] = 4'hE;
    Number7[14][7] = 4'hC;
    Number7[15][7] = 4'hC;
    Number7[16][7] = 4'hC;
    Number7[17][7] = 4'hC;
    Number7[18][7] = 4'hC;
    Number7[19][7] = 4'hD;
    Number7[20][7] = 4'hF;
    Number7[21][7] = 4'hF;
    Number7[22][7] = 4'hF;
    Number7[0][8] = 4'hF;
    Number7[1][8] = 4'hF;
    Number7[2][8] = 4'hF;
    Number7[3][8] = 4'hF;
    Number7[4][8] = 4'hF;
    Number7[5][8] = 4'hF;
    Number7[6][8] = 4'hF;
    Number7[7][8] = 4'hF;
    Number7[8][8] = 4'hF;
    Number7[9][8] = 4'hF;
    Number7[10][8] = 4'hF;
    Number7[11][8] = 4'hF;
    Number7[12][8] = 4'hF;
    Number7[13][8] = 4'hD;
    Number7[14][8] = 4'hC;
    Number7[15][8] = 4'hC;
    Number7[16][8] = 4'hC;
    Number7[17][8] = 4'hC;
    Number7[18][8] = 4'hC;
    Number7[19][8] = 4'hF;
    Number7[20][8] = 4'hF;
    Number7[21][8] = 4'hF;
    Number7[22][8] = 4'hF;
    Number7[0][9] = 4'hF;
    Number7[1][9] = 4'hF;
    Number7[2][9] = 4'hF;
    Number7[3][9] = 4'hF;
    Number7[4][9] = 4'hF;
    Number7[5][9] = 4'hF;
    Number7[6][9] = 4'hF;
    Number7[7][9] = 4'hF;
    Number7[8][9] = 4'hF;
    Number7[9][9] = 4'hF;
    Number7[10][9] = 4'hF;
    Number7[11][9] = 4'hF;
    Number7[12][9] = 4'hE;
    Number7[13][9] = 4'hC;
    Number7[14][9] = 4'hC;
    Number7[15][9] = 4'hC;
    Number7[16][9] = 4'hC;
    Number7[17][9] = 4'hC;
    Number7[18][9] = 4'hD;
    Number7[19][9] = 4'hF;
    Number7[20][9] = 4'hF;
    Number7[21][9] = 4'hF;
    Number7[22][9] = 4'hF;
    Number7[0][10] = 4'hF;
    Number7[1][10] = 4'hF;
    Number7[2][10] = 4'hF;
    Number7[3][10] = 4'hF;
    Number7[4][10] = 4'hF;
    Number7[5][10] = 4'hF;
    Number7[6][10] = 4'hF;
    Number7[7][10] = 4'hF;
    Number7[8][10] = 4'hF;
    Number7[9][10] = 4'hF;
    Number7[10][10] = 4'hF;
    Number7[11][10] = 4'hF;
    Number7[12][10] = 4'hD;
    Number7[13][10] = 4'hC;
    Number7[14][10] = 4'hC;
    Number7[15][10] = 4'hC;
    Number7[16][10] = 4'hC;
    Number7[17][10] = 4'hC;
    Number7[18][10] = 4'hF;
    Number7[19][10] = 4'hF;
    Number7[20][10] = 4'hF;
    Number7[21][10] = 4'hF;
    Number7[22][10] = 4'hF;
    Number7[0][11] = 4'hF;
    Number7[1][11] = 4'hF;
    Number7[2][11] = 4'hF;
    Number7[3][11] = 4'hF;
    Number7[4][11] = 4'hF;
    Number7[5][11] = 4'hF;
    Number7[6][11] = 4'hF;
    Number7[7][11] = 4'hF;
    Number7[8][11] = 4'hF;
    Number7[9][11] = 4'hF;
    Number7[10][11] = 4'hF;
    Number7[11][11] = 4'hF;
    Number7[12][11] = 4'hC;
    Number7[13][11] = 4'hC;
    Number7[14][11] = 4'hC;
    Number7[15][11] = 4'hC;
    Number7[16][11] = 4'hC;
    Number7[17][11] = 4'hD;
    Number7[18][11] = 4'hF;
    Number7[19][11] = 4'hF;
    Number7[20][11] = 4'hF;
    Number7[21][11] = 4'hF;
    Number7[22][11] = 4'hF;
    Number7[0][12] = 4'hF;
    Number7[1][12] = 4'hF;
    Number7[2][12] = 4'hF;
    Number7[3][12] = 4'hF;
    Number7[4][12] = 4'hF;
    Number7[5][12] = 4'hF;
    Number7[6][12] = 4'hF;
    Number7[7][12] = 4'hF;
    Number7[8][12] = 4'hF;
    Number7[9][12] = 4'hF;
    Number7[10][12] = 4'hF;
    Number7[11][12] = 4'hD;
    Number7[12][12] = 4'hC;
    Number7[13][12] = 4'hC;
    Number7[14][12] = 4'hC;
    Number7[15][12] = 4'hC;
    Number7[16][12] = 4'hC;
    Number7[17][12] = 4'hE;
    Number7[18][12] = 4'hF;
    Number7[19][12] = 4'hF;
    Number7[20][12] = 4'hF;
    Number7[21][12] = 4'hF;
    Number7[22][12] = 4'hF;
    Number7[0][13] = 4'hF;
    Number7[1][13] = 4'hF;
    Number7[2][13] = 4'hF;
    Number7[3][13] = 4'hF;
    Number7[4][13] = 4'hF;
    Number7[5][13] = 4'hF;
    Number7[6][13] = 4'hF;
    Number7[7][13] = 4'hF;
    Number7[8][13] = 4'hF;
    Number7[9][13] = 4'hF;
    Number7[10][13] = 4'hF;
    Number7[11][13] = 4'hC;
    Number7[12][13] = 4'hC;
    Number7[13][13] = 4'hC;
    Number7[14][13] = 4'hC;
    Number7[15][13] = 4'hC;
    Number7[16][13] = 4'hD;
    Number7[17][13] = 4'hF;
    Number7[18][13] = 4'hF;
    Number7[19][13] = 4'hF;
    Number7[20][13] = 4'hF;
    Number7[21][13] = 4'hF;
    Number7[22][13] = 4'hF;
    Number7[0][14] = 4'hF;
    Number7[1][14] = 4'hF;
    Number7[2][14] = 4'hF;
    Number7[3][14] = 4'hF;
    Number7[4][14] = 4'hF;
    Number7[5][14] = 4'hF;
    Number7[6][14] = 4'hF;
    Number7[7][14] = 4'hF;
    Number7[8][14] = 4'hF;
    Number7[9][14] = 4'hF;
    Number7[10][14] = 4'hD;
    Number7[11][14] = 4'hC;
    Number7[12][14] = 4'hC;
    Number7[13][14] = 4'hC;
    Number7[14][14] = 4'hC;
    Number7[15][14] = 4'hC;
    Number7[16][14] = 4'hD;
    Number7[17][14] = 4'hF;
    Number7[18][14] = 4'hF;
    Number7[19][14] = 4'hF;
    Number7[20][14] = 4'hF;
    Number7[21][14] = 4'hF;
    Number7[22][14] = 4'hF;
    Number7[0][15] = 4'hF;
    Number7[1][15] = 4'hF;
    Number7[2][15] = 4'hF;
    Number7[3][15] = 4'hF;
    Number7[4][15] = 4'hF;
    Number7[5][15] = 4'hF;
    Number7[6][15] = 4'hF;
    Number7[7][15] = 4'hF;
    Number7[8][15] = 4'hF;
    Number7[9][15] = 4'hF;
    Number7[10][15] = 4'hC;
    Number7[11][15] = 4'hC;
    Number7[12][15] = 4'hC;
    Number7[13][15] = 4'hC;
    Number7[14][15] = 4'hC;
    Number7[15][15] = 4'hC;
    Number7[16][15] = 4'hF;
    Number7[17][15] = 4'hF;
    Number7[18][15] = 4'hF;
    Number7[19][15] = 4'hF;
    Number7[20][15] = 4'hF;
    Number7[21][15] = 4'hF;
    Number7[22][15] = 4'hF;
    Number7[0][16] = 4'hF;
    Number7[1][16] = 4'hF;
    Number7[2][16] = 4'hF;
    Number7[3][16] = 4'hF;
    Number7[4][16] = 4'hF;
    Number7[5][16] = 4'hF;
    Number7[6][16] = 4'hF;
    Number7[7][16] = 4'hF;
    Number7[8][16] = 4'hF;
    Number7[9][16] = 4'hE;
    Number7[10][16] = 4'hC;
    Number7[11][16] = 4'hC;
    Number7[12][16] = 4'hC;
    Number7[13][16] = 4'hC;
    Number7[14][16] = 4'hC;
    Number7[15][16] = 4'hD;
    Number7[16][16] = 4'hF;
    Number7[17][16] = 4'hF;
    Number7[18][16] = 4'hF;
    Number7[19][16] = 4'hF;
    Number7[20][16] = 4'hF;
    Number7[21][16] = 4'hF;
    Number7[22][16] = 4'hF;
    Number7[0][17] = 4'hF;
    Number7[1][17] = 4'hF;
    Number7[2][17] = 4'hF;
    Number7[3][17] = 4'hF;
    Number7[4][17] = 4'hF;
    Number7[5][17] = 4'hF;
    Number7[6][17] = 4'hF;
    Number7[7][17] = 4'hF;
    Number7[8][17] = 4'hF;
    Number7[9][17] = 4'hD;
    Number7[10][17] = 4'hC;
    Number7[11][17] = 4'hC;
    Number7[12][17] = 4'hC;
    Number7[13][17] = 4'hC;
    Number7[14][17] = 4'hC;
    Number7[15][17] = 4'hF;
    Number7[16][17] = 4'hF;
    Number7[17][17] = 4'hF;
    Number7[18][17] = 4'hF;
    Number7[19][17] = 4'hF;
    Number7[20][17] = 4'hF;
    Number7[21][17] = 4'hF;
    Number7[22][17] = 4'hF;
    Number7[0][18] = 4'hF;
    Number7[1][18] = 4'hF;
    Number7[2][18] = 4'hF;
    Number7[3][18] = 4'hF;
    Number7[4][18] = 4'hF;
    Number7[5][18] = 4'hF;
    Number7[6][18] = 4'hF;
    Number7[7][18] = 4'hF;
    Number7[8][18] = 4'hE;
    Number7[9][18] = 4'hC;
    Number7[10][18] = 4'hC;
    Number7[11][18] = 4'hC;
    Number7[12][18] = 4'hC;
    Number7[13][18] = 4'hC;
    Number7[14][18] = 4'hD;
    Number7[15][18] = 4'hF;
    Number7[16][18] = 4'hF;
    Number7[17][18] = 4'hF;
    Number7[18][18] = 4'hF;
    Number7[19][18] = 4'hF;
    Number7[20][18] = 4'hF;
    Number7[21][18] = 4'hF;
    Number7[22][18] = 4'hF;
    Number7[0][19] = 4'hF;
    Number7[1][19] = 4'hF;
    Number7[2][19] = 4'hF;
    Number7[3][19] = 4'hF;
    Number7[4][19] = 4'hF;
    Number7[5][19] = 4'hF;
    Number7[6][19] = 4'hF;
    Number7[7][19] = 4'hF;
    Number7[8][19] = 4'hD;
    Number7[9][19] = 4'hC;
    Number7[10][19] = 4'hC;
    Number7[11][19] = 4'hC;
    Number7[12][19] = 4'hC;
    Number7[13][19] = 4'hC;
    Number7[14][19] = 4'hE;
    Number7[15][19] = 4'hF;
    Number7[16][19] = 4'hF;
    Number7[17][19] = 4'hF;
    Number7[18][19] = 4'hF;
    Number7[19][19] = 4'hF;
    Number7[20][19] = 4'hF;
    Number7[21][19] = 4'hF;
    Number7[22][19] = 4'hF;
    Number7[0][20] = 4'hF;
    Number7[1][20] = 4'hF;
    Number7[2][20] = 4'hF;
    Number7[3][20] = 4'hF;
    Number7[4][20] = 4'hF;
    Number7[5][20] = 4'hF;
    Number7[6][20] = 4'hF;
    Number7[7][20] = 4'hE;
    Number7[8][20] = 4'hC;
    Number7[9][20] = 4'hC;
    Number7[10][20] = 4'hC;
    Number7[11][20] = 4'hC;
    Number7[12][20] = 4'hC;
    Number7[13][20] = 4'hD;
    Number7[14][20] = 4'hF;
    Number7[15][20] = 4'hF;
    Number7[16][20] = 4'hF;
    Number7[17][20] = 4'hF;
    Number7[18][20] = 4'hF;
    Number7[19][20] = 4'hF;
    Number7[20][20] = 4'hF;
    Number7[21][20] = 4'hF;
    Number7[22][20] = 4'hF;
    Number7[0][21] = 4'hF;
    Number7[1][21] = 4'hF;
    Number7[2][21] = 4'hF;
    Number7[3][21] = 4'hF;
    Number7[4][21] = 4'hF;
    Number7[5][21] = 4'hF;
    Number7[6][21] = 4'hF;
    Number7[7][21] = 4'hD;
    Number7[8][21] = 4'hC;
    Number7[9][21] = 4'hC;
    Number7[10][21] = 4'hC;
    Number7[11][21] = 4'hC;
    Number7[12][21] = 4'hC;
    Number7[13][21] = 4'hD;
    Number7[14][21] = 4'hF;
    Number7[15][21] = 4'hF;
    Number7[16][21] = 4'hF;
    Number7[17][21] = 4'hF;
    Number7[18][21] = 4'hF;
    Number7[19][21] = 4'hF;
    Number7[20][21] = 4'hF;
    Number7[21][21] = 4'hF;
    Number7[22][21] = 4'hF;
    Number7[0][22] = 4'hF;
    Number7[1][22] = 4'hF;
    Number7[2][22] = 4'hF;
    Number7[3][22] = 4'hF;
    Number7[4][22] = 4'hF;
    Number7[5][22] = 4'hF;
    Number7[6][22] = 4'hF;
    Number7[7][22] = 4'hC;
    Number7[8][22] = 4'hC;
    Number7[9][22] = 4'hC;
    Number7[10][22] = 4'hC;
    Number7[11][22] = 4'hC;
    Number7[12][22] = 4'hC;
    Number7[13][22] = 4'hF;
    Number7[14][22] = 4'hF;
    Number7[15][22] = 4'hF;
    Number7[16][22] = 4'hF;
    Number7[17][22] = 4'hF;
    Number7[18][22] = 4'hF;
    Number7[19][22] = 4'hF;
    Number7[20][22] = 4'hF;
    Number7[21][22] = 4'hF;
    Number7[22][22] = 4'hF;
    Number7[0][23] = 4'hF;
    Number7[1][23] = 4'hF;
    Number7[2][23] = 4'hF;
    Number7[3][23] = 4'hF;
    Number7[4][23] = 4'hF;
    Number7[5][23] = 4'hF;
    Number7[6][23] = 4'hD;
    Number7[7][23] = 4'hC;
    Number7[8][23] = 4'hC;
    Number7[9][23] = 4'hC;
    Number7[10][23] = 4'hC;
    Number7[11][23] = 4'hC;
    Number7[12][23] = 4'hD;
    Number7[13][23] = 4'hF;
    Number7[14][23] = 4'hF;
    Number7[15][23] = 4'hF;
    Number7[16][23] = 4'hF;
    Number7[17][23] = 4'hF;
    Number7[18][23] = 4'hF;
    Number7[19][23] = 4'hF;
    Number7[20][23] = 4'hF;
    Number7[21][23] = 4'hF;
    Number7[22][23] = 4'hF;
    Number7[0][24] = 4'hF;
    Number7[1][24] = 4'hF;
    Number7[2][24] = 4'hF;
    Number7[3][24] = 4'hF;
    Number7[4][24] = 4'hF;
    Number7[5][24] = 4'hF;
    Number7[6][24] = 4'hC;
    Number7[7][24] = 4'hC;
    Number7[8][24] = 4'hC;
    Number7[9][24] = 4'hC;
    Number7[10][24] = 4'hC;
    Number7[11][24] = 4'hC;
    Number7[12][24] = 4'hF;
    Number7[13][24] = 4'hF;
    Number7[14][24] = 4'hF;
    Number7[15][24] = 4'hF;
    Number7[16][24] = 4'hF;
    Number7[17][24] = 4'hF;
    Number7[18][24] = 4'hF;
    Number7[19][24] = 4'hF;
    Number7[20][24] = 4'hF;
    Number7[21][24] = 4'hF;
    Number7[22][24] = 4'hF;
    Number7[0][25] = 4'hF;
    Number7[1][25] = 4'hF;
    Number7[2][25] = 4'hF;
    Number7[3][25] = 4'hF;
    Number7[4][25] = 4'hF;
    Number7[5][25] = 4'hD;
    Number7[6][25] = 4'hC;
    Number7[7][25] = 4'hC;
    Number7[8][25] = 4'hC;
    Number7[9][25] = 4'hC;
    Number7[10][25] = 4'hC;
    Number7[11][25] = 4'hD;
    Number7[12][25] = 4'hF;
    Number7[13][25] = 4'hF;
    Number7[14][25] = 4'hF;
    Number7[15][25] = 4'hF;
    Number7[16][25] = 4'hF;
    Number7[17][25] = 4'hF;
    Number7[18][25] = 4'hF;
    Number7[19][25] = 4'hF;
    Number7[20][25] = 4'hF;
    Number7[21][25] = 4'hF;
    Number7[22][25] = 4'hF;
    Number7[0][26] = 4'hF;
    Number7[1][26] = 4'hF;
    Number7[2][26] = 4'hF;
    Number7[3][26] = 4'hF;
    Number7[4][26] = 4'hF;
    Number7[5][26] = 4'hD;
    Number7[6][26] = 4'hC;
    Number7[7][26] = 4'hC;
    Number7[8][26] = 4'hC;
    Number7[9][26] = 4'hC;
    Number7[10][26] = 4'hC;
    Number7[11][26] = 4'hE;
    Number7[12][26] = 4'hF;
    Number7[13][26] = 4'hF;
    Number7[14][26] = 4'hF;
    Number7[15][26] = 4'hF;
    Number7[16][26] = 4'hF;
    Number7[17][26] = 4'hF;
    Number7[18][26] = 4'hF;
    Number7[19][26] = 4'hF;
    Number7[20][26] = 4'hF;
    Number7[21][26] = 4'hF;
    Number7[22][26] = 4'hF;
    Number7[0][27] = 4'hF;
    Number7[1][27] = 4'hF;
    Number7[2][27] = 4'hF;
    Number7[3][27] = 4'hF;
    Number7[4][27] = 4'hF;
    Number7[5][27] = 4'hF;
    Number7[6][27] = 4'hF;
    Number7[7][27] = 4'hF;
    Number7[8][27] = 4'hF;
    Number7[9][27] = 4'hF;
    Number7[10][27] = 4'hF;
    Number7[11][27] = 4'hF;
    Number7[12][27] = 4'hF;
    Number7[13][27] = 4'hF;
    Number7[14][27] = 4'hF;
    Number7[15][27] = 4'hF;
    Number7[16][27] = 4'hF;
    Number7[17][27] = 4'hF;
    Number7[18][27] = 4'hF;
    Number7[19][27] = 4'hF;
    Number7[20][27] = 4'hF;
    Number7[21][27] = 4'hF;
    Number7[22][27] = 4'hF;
    Number7[0][28] = 4'hF;
    Number7[1][28] = 4'hF;
    Number7[2][28] = 4'hF;
    Number7[3][28] = 4'hF;
    Number7[4][28] = 4'hF;
    Number7[5][28] = 4'hF;
    Number7[6][28] = 4'hF;
    Number7[7][28] = 4'hF;
    Number7[8][28] = 4'hF;
    Number7[9][28] = 4'hF;
    Number7[10][28] = 4'hF;
    Number7[11][28] = 4'hF;
    Number7[12][28] = 4'hF;
    Number7[13][28] = 4'hF;
    Number7[14][28] = 4'hF;
    Number7[15][28] = 4'hF;
    Number7[16][28] = 4'hF;
    Number7[17][28] = 4'hF;
    Number7[18][28] = 4'hF;
    Number7[19][28] = 4'hF;
    Number7[20][28] = 4'hF;
    Number7[21][28] = 4'hF;
    Number7[22][28] = 4'hF;

// Number 8
    Number8[0][0] = 4'hF;
    Number8[1][0] = 4'hF;
    Number8[2][0] = 4'hF;
    Number8[3][0] = 4'hF;
    Number8[4][0] = 4'hF;
    Number8[5][0] = 4'hF;
    Number8[6][0] = 4'hF;
    Number8[7][0] = 4'hF;
    Number8[8][0] = 4'hF;
    Number8[9][0] = 4'hF;
    Number8[10][0] = 4'hF;
    Number8[11][0] = 4'hF;
    Number8[12][0] = 4'hF;
    Number8[13][0] = 4'hF;
    Number8[14][0] = 4'hF;
    Number8[15][0] = 4'hF;
    Number8[16][0] = 4'hF;
    Number8[17][0] = 4'hF;
    Number8[18][0] = 4'hF;
    Number8[19][0] = 4'hF;
    Number8[20][0] = 4'hF;
    Number8[21][0] = 4'hF;
    Number8[22][0] = 4'hF;
    Number8[0][1] = 4'hF;
    Number8[1][1] = 4'hF;
    Number8[2][1] = 4'hF;
    Number8[3][1] = 4'hF;
    Number8[4][1] = 4'hF;
    Number8[5][1] = 4'hF;
    Number8[6][1] = 4'hF;
    Number8[7][1] = 4'hF;
    Number8[8][1] = 4'hF;
    Number8[9][1] = 4'hF;
    Number8[10][1] = 4'hF;
    Number8[11][1] = 4'hF;
    Number8[12][1] = 4'hF;
    Number8[13][1] = 4'hF;
    Number8[14][1] = 4'hF;
    Number8[15][1] = 4'hF;
    Number8[16][1] = 4'hF;
    Number8[17][1] = 4'hF;
    Number8[18][1] = 4'hF;
    Number8[19][1] = 4'hF;
    Number8[20][1] = 4'hF;
    Number8[21][1] = 4'hF;
    Number8[22][1] = 4'hF;
    Number8[0][2] = 4'hF;
    Number8[1][2] = 4'hF;
    Number8[2][2] = 4'hF;
    Number8[3][2] = 4'hF;
    Number8[4][2] = 4'hF;
    Number8[5][2] = 4'hF;
    Number8[6][2] = 4'hF;
    Number8[7][2] = 4'hD;
    Number8[8][2] = 4'hD;
    Number8[9][2] = 4'hC;
    Number8[10][2] = 4'hC;
    Number8[11][2] = 4'hC;
    Number8[12][2] = 4'hC;
    Number8[13][2] = 4'hC;
    Number8[14][2] = 4'hC;
    Number8[15][2] = 4'hD;
    Number8[16][2] = 4'hE;
    Number8[17][2] = 4'hF;
    Number8[18][2] = 4'hF;
    Number8[19][2] = 4'hF;
    Number8[20][2] = 4'hF;
    Number8[21][2] = 4'hF;
    Number8[22][2] = 4'hF;
    Number8[0][3] = 4'hF;
    Number8[1][3] = 4'hF;
    Number8[2][3] = 4'hF;
    Number8[3][3] = 4'hF;
    Number8[4][3] = 4'hF;
    Number8[5][3] = 4'hE;
    Number8[6][3] = 4'hC;
    Number8[7][3] = 4'hC;
    Number8[8][3] = 4'hC;
    Number8[9][3] = 4'hC;
    Number8[10][3] = 4'hC;
    Number8[11][3] = 4'hC;
    Number8[12][3] = 4'hC;
    Number8[13][3] = 4'hC;
    Number8[14][3] = 4'hC;
    Number8[15][3] = 4'hC;
    Number8[16][3] = 4'hC;
    Number8[17][3] = 4'hD;
    Number8[18][3] = 4'hF;
    Number8[19][3] = 4'hF;
    Number8[20][3] = 4'hF;
    Number8[21][3] = 4'hF;
    Number8[22][3] = 4'hF;
    Number8[0][4] = 4'hF;
    Number8[1][4] = 4'hF;
    Number8[2][4] = 4'hF;
    Number8[3][4] = 4'hF;
    Number8[4][4] = 4'hE;
    Number8[5][4] = 4'hC;
    Number8[6][4] = 4'hC;
    Number8[7][4] = 4'hC;
    Number8[8][4] = 4'hC;
    Number8[9][4] = 4'hC;
    Number8[10][4] = 4'hC;
    Number8[11][4] = 4'hC;
    Number8[12][4] = 4'hC;
    Number8[13][4] = 4'hC;
    Number8[14][4] = 4'hC;
    Number8[15][4] = 4'hC;
    Number8[16][4] = 4'hC;
    Number8[17][4] = 4'hC;
    Number8[18][4] = 4'hC;
    Number8[19][4] = 4'hF;
    Number8[20][4] = 4'hF;
    Number8[21][4] = 4'hF;
    Number8[22][4] = 4'hF;
    Number8[0][5] = 4'hF;
    Number8[1][5] = 4'hF;
    Number8[2][5] = 4'hF;
    Number8[3][5] = 4'hF;
    Number8[4][5] = 4'hC;
    Number8[5][5] = 4'hC;
    Number8[6][5] = 4'hC;
    Number8[7][5] = 4'hC;
    Number8[8][5] = 4'hC;
    Number8[9][5] = 4'hC;
    Number8[10][5] = 4'hC;
    Number8[11][5] = 4'hC;
    Number8[12][5] = 4'hC;
    Number8[13][5] = 4'hC;
    Number8[14][5] = 4'hC;
    Number8[15][5] = 4'hC;
    Number8[16][5] = 4'hC;
    Number8[17][5] = 4'hC;
    Number8[18][5] = 4'hC;
    Number8[19][5] = 4'hD;
    Number8[20][5] = 4'hF;
    Number8[21][5] = 4'hF;
    Number8[22][5] = 4'hF;
    Number8[0][6] = 4'hF;
    Number8[1][6] = 4'hF;
    Number8[2][6] = 4'hF;
    Number8[3][6] = 4'hD;
    Number8[4][6] = 4'hC;
    Number8[5][6] = 4'hC;
    Number8[6][6] = 4'hC;
    Number8[7][6] = 4'hC;
    Number8[8][6] = 4'hC;
    Number8[9][6] = 4'hD;
    Number8[10][6] = 4'hE;
    Number8[11][6] = 4'hF;
    Number8[12][6] = 4'hE;
    Number8[13][6] = 4'hD;
    Number8[14][6] = 4'hC;
    Number8[15][6] = 4'hC;
    Number8[16][6] = 4'hC;
    Number8[17][6] = 4'hC;
    Number8[18][6] = 4'hC;
    Number8[19][6] = 4'hD;
    Number8[20][6] = 4'hF;
    Number8[21][6] = 4'hF;
    Number8[22][6] = 4'hF;
    Number8[0][7] = 4'hF;
    Number8[1][7] = 4'hF;
    Number8[2][7] = 4'hF;
    Number8[3][7] = 4'hD;
    Number8[4][7] = 4'hC;
    Number8[5][7] = 4'hC;
    Number8[6][7] = 4'hC;
    Number8[7][7] = 4'hC;
    Number8[8][7] = 4'hD;
    Number8[9][7] = 4'hF;
    Number8[10][7] = 4'hF;
    Number8[11][7] = 4'hF;
    Number8[12][7] = 4'hF;
    Number8[13][7] = 4'hF;
    Number8[14][7] = 4'hD;
    Number8[15][7] = 4'hC;
    Number8[16][7] = 4'hC;
    Number8[17][7] = 4'hC;
    Number8[18][7] = 4'hC;
    Number8[19][7] = 4'hC;
    Number8[20][7] = 4'hF;
    Number8[21][7] = 4'hF;
    Number8[22][7] = 4'hF;
    Number8[0][8] = 4'hF;
    Number8[1][8] = 4'hF;
    Number8[2][8] = 4'hF;
    Number8[3][8] = 4'hD;
    Number8[4][8] = 4'hC;
    Number8[5][8] = 4'hC;
    Number8[6][8] = 4'hC;
    Number8[7][8] = 4'hC;
    Number8[8][8] = 4'hD;
    Number8[9][8] = 4'hF;
    Number8[10][8] = 4'hF;
    Number8[11][8] = 4'hF;
    Number8[12][8] = 4'hF;
    Number8[13][8] = 4'hF;
    Number8[14][8] = 4'hE;
    Number8[15][8] = 4'hC;
    Number8[16][8] = 4'hC;
    Number8[17][8] = 4'hC;
    Number8[18][8] = 4'hC;
    Number8[19][8] = 4'hC;
    Number8[20][8] = 4'hF;
    Number8[21][8] = 4'hF;
    Number8[22][8] = 4'hF;
    Number8[0][9] = 4'hF;
    Number8[1][9] = 4'hF;
    Number8[2][9] = 4'hF;
    Number8[3][9] = 4'hD;
    Number8[4][9] = 4'hC;
    Number8[5][9] = 4'hC;
    Number8[6][9] = 4'hC;
    Number8[7][9] = 4'hC;
    Number8[8][9] = 4'hD;
    Number8[9][9] = 4'hF;
    Number8[10][9] = 4'hF;
    Number8[11][9] = 4'hF;
    Number8[12][9] = 4'hF;
    Number8[13][9] = 4'hF;
    Number8[14][9] = 4'hD;
    Number8[15][9] = 4'hC;
    Number8[16][9] = 4'hC;
    Number8[17][9] = 4'hC;
    Number8[18][9] = 4'hC;
    Number8[19][9] = 4'hD;
    Number8[20][9] = 4'hF;
    Number8[21][9] = 4'hF;
    Number8[22][9] = 4'hF;
    Number8[0][10] = 4'hF;
    Number8[1][10] = 4'hF;
    Number8[2][10] = 4'hF;
    Number8[3][10] = 4'hE;
    Number8[4][10] = 4'hC;
    Number8[5][10] = 4'hC;
    Number8[6][10] = 4'hC;
    Number8[7][10] = 4'hC;
    Number8[8][10] = 4'hC;
    Number8[9][10] = 4'hD;
    Number8[10][10] = 4'hF;
    Number8[11][10] = 4'hF;
    Number8[12][10] = 4'hF;
    Number8[13][10] = 4'hE;
    Number8[14][10] = 4'hC;
    Number8[15][10] = 4'hC;
    Number8[16][10] = 4'hC;
    Number8[17][10] = 4'hC;
    Number8[18][10] = 4'hC;
    Number8[19][10] = 4'hE;
    Number8[20][10] = 4'hF;
    Number8[21][10] = 4'hF;
    Number8[22][10] = 4'hF;
    Number8[0][11] = 4'hF;
    Number8[1][11] = 4'hF;
    Number8[2][11] = 4'hF;
    Number8[3][11] = 4'hF;
    Number8[4][11] = 4'hC;
    Number8[5][11] = 4'hC;
    Number8[6][11] = 4'hC;
    Number8[7][11] = 4'hC;
    Number8[8][11] = 4'hC;
    Number8[9][11] = 4'hC;
    Number8[10][11] = 4'hD;
    Number8[11][11] = 4'hE;
    Number8[12][11] = 4'hE;
    Number8[13][11] = 4'hC;
    Number8[14][11] = 4'hC;
    Number8[15][11] = 4'hC;
    Number8[16][11] = 4'hC;
    Number8[17][11] = 4'hC;
    Number8[18][11] = 4'hD;
    Number8[19][11] = 4'hF;
    Number8[20][11] = 4'hF;
    Number8[21][11] = 4'hF;
    Number8[22][11] = 4'hF;
    Number8[0][12] = 4'hF;
    Number8[1][12] = 4'hF;
    Number8[2][12] = 4'hF;
    Number8[3][12] = 4'hF;
    Number8[4][12] = 4'hE;
    Number8[5][12] = 4'hC;
    Number8[6][12] = 4'hC;
    Number8[7][12] = 4'hC;
    Number8[8][12] = 4'hC;
    Number8[9][12] = 4'hC;
    Number8[10][12] = 4'hC;
    Number8[11][12] = 4'hC;
    Number8[12][12] = 4'hC;
    Number8[13][12] = 4'hC;
    Number8[14][12] = 4'hC;
    Number8[15][12] = 4'hC;
    Number8[16][12] = 4'hC;
    Number8[17][12] = 4'hD;
    Number8[18][12] = 4'hF;
    Number8[19][12] = 4'hF;
    Number8[20][12] = 4'hF;
    Number8[21][12] = 4'hF;
    Number8[22][12] = 4'hF;
    Number8[0][13] = 4'hF;
    Number8[1][13] = 4'hF;
    Number8[2][13] = 4'hF;
    Number8[3][13] = 4'hF;
    Number8[4][13] = 4'hF;
    Number8[5][13] = 4'hE;
    Number8[6][13] = 4'hD;
    Number8[7][13] = 4'hC;
    Number8[8][13] = 4'hC;
    Number8[9][13] = 4'hC;
    Number8[10][13] = 4'hC;
    Number8[11][13] = 4'hC;
    Number8[12][13] = 4'hC;
    Number8[13][13] = 4'hC;
    Number8[14][13] = 4'hC;
    Number8[15][13] = 4'hC;
    Number8[16][13] = 4'hE;
    Number8[17][13] = 4'hF;
    Number8[18][13] = 4'hF;
    Number8[19][13] = 4'hF;
    Number8[20][13] = 4'hF;
    Number8[21][13] = 4'hF;
    Number8[22][13] = 4'hF;
    Number8[0][14] = 4'hF;
    Number8[1][14] = 4'hF;
    Number8[2][14] = 4'hF;
    Number8[3][14] = 4'hF;
    Number8[4][14] = 4'hF;
    Number8[5][14] = 4'hF;
    Number8[6][14] = 4'hF;
    Number8[7][14] = 4'hD;
    Number8[8][14] = 4'hC;
    Number8[9][14] = 4'hC;
    Number8[10][14] = 4'hC;
    Number8[11][14] = 4'hC;
    Number8[12][14] = 4'hC;
    Number8[13][14] = 4'hC;
    Number8[14][14] = 4'hC;
    Number8[15][14] = 4'hC;
    Number8[16][14] = 4'hD;
    Number8[17][14] = 4'hE;
    Number8[18][14] = 4'hF;
    Number8[19][14] = 4'hF;
    Number8[20][14] = 4'hF;
    Number8[21][14] = 4'hF;
    Number8[22][14] = 4'hF;
    Number8[0][15] = 4'hF;
    Number8[1][15] = 4'hF;
    Number8[2][15] = 4'hF;
    Number8[3][15] = 4'hF;
    Number8[4][15] = 4'hF;
    Number8[5][15] = 4'hD;
    Number8[6][15] = 4'hC;
    Number8[7][15] = 4'hC;
    Number8[8][15] = 4'hC;
    Number8[9][15] = 4'hC;
    Number8[10][15] = 4'hC;
    Number8[11][15] = 4'hC;
    Number8[12][15] = 4'hC;
    Number8[13][15] = 4'hC;
    Number8[14][15] = 4'hC;
    Number8[15][15] = 4'hC;
    Number8[16][15] = 4'hC;
    Number8[17][15] = 4'hC;
    Number8[18][15] = 4'hE;
    Number8[19][15] = 4'hF;
    Number8[20][15] = 4'hF;
    Number8[21][15] = 4'hF;
    Number8[22][15] = 4'hF;
    Number8[0][16] = 4'hF;
    Number8[1][16] = 4'hF;
    Number8[2][16] = 4'hF;
    Number8[3][16] = 4'hF;
    Number8[4][16] = 4'hD;
    Number8[5][16] = 4'hC;
    Number8[6][16] = 4'hC;
    Number8[7][16] = 4'hC;
    Number8[8][16] = 4'hC;
    Number8[9][16] = 4'hC;
    Number8[10][16] = 4'hD;
    Number8[11][16] = 4'hD;
    Number8[12][16] = 4'hC;
    Number8[13][16] = 4'hC;
    Number8[14][16] = 4'hC;
    Number8[15][16] = 4'hC;
    Number8[16][16] = 4'hC;
    Number8[17][16] = 4'hC;
    Number8[18][16] = 4'hC;
    Number8[19][16] = 4'hE;
    Number8[20][16] = 4'hF;
    Number8[21][16] = 4'hF;
    Number8[22][16] = 4'hF;
    Number8[0][17] = 4'hF;
    Number8[1][17] = 4'hF;
    Number8[2][17] = 4'hF;
    Number8[3][17] = 4'hD;
    Number8[4][17] = 4'hC;
    Number8[5][17] = 4'hC;
    Number8[6][17] = 4'hC;
    Number8[7][17] = 4'hC;
    Number8[8][17] = 4'hC;
    Number8[9][17] = 4'hD;
    Number8[10][17] = 4'hF;
    Number8[11][17] = 4'hF;
    Number8[12][17] = 4'hF;
    Number8[13][17] = 4'hD;
    Number8[14][17] = 4'hC;
    Number8[15][17] = 4'hC;
    Number8[16][17] = 4'hC;
    Number8[17][17] = 4'hC;
    Number8[18][17] = 4'hC;
    Number8[19][17] = 4'hC;
    Number8[20][17] = 4'hF;
    Number8[21][17] = 4'hF;
    Number8[22][17] = 4'hF;
    Number8[0][18] = 4'hF;
    Number8[1][18] = 4'hF;
    Number8[2][18] = 4'hF;
    Number8[3][18] = 4'hC;
    Number8[4][18] = 4'hC;
    Number8[5][18] = 4'hC;
    Number8[6][18] = 4'hC;
    Number8[7][18] = 4'hC;
    Number8[8][18] = 4'hD;
    Number8[9][18] = 4'hF;
    Number8[10][18] = 4'hF;
    Number8[11][18] = 4'hF;
    Number8[12][18] = 4'hF;
    Number8[13][18] = 4'hF;
    Number8[14][18] = 4'hE;
    Number8[15][18] = 4'hC;
    Number8[16][18] = 4'hC;
    Number8[17][18] = 4'hC;
    Number8[18][18] = 4'hC;
    Number8[19][18] = 4'hC;
    Number8[20][18] = 4'hD;
    Number8[21][18] = 4'hF;
    Number8[22][18] = 4'hF;
    Number8[0][19] = 4'hF;
    Number8[1][19] = 4'hF;
    Number8[2][19] = 4'hE;
    Number8[3][19] = 4'hC;
    Number8[4][19] = 4'hC;
    Number8[5][19] = 4'hC;
    Number8[6][19] = 4'hC;
    Number8[7][19] = 4'hC;
    Number8[8][19] = 4'hF;
    Number8[9][19] = 4'hF;
    Number8[10][19] = 4'hF;
    Number8[11][19] = 4'hF;
    Number8[12][19] = 4'hF;
    Number8[13][19] = 4'hF;
    Number8[14][19] = 4'hF;
    Number8[15][19] = 4'hD;
    Number8[16][19] = 4'hC;
    Number8[17][19] = 4'hC;
    Number8[18][19] = 4'hC;
    Number8[19][19] = 4'hC;
    Number8[20][19] = 4'hD;
    Number8[21][19] = 4'hF;
    Number8[22][19] = 4'hF;
    Number8[0][20] = 4'hF;
    Number8[1][20] = 4'hF;
    Number8[2][20] = 4'hD;
    Number8[3][20] = 4'hC;
    Number8[4][20] = 4'hC;
    Number8[5][20] = 4'hC;
    Number8[6][20] = 4'hC;
    Number8[7][20] = 4'hC;
    Number8[8][20] = 4'hF;
    Number8[9][20] = 4'hF;
    Number8[10][20] = 4'hF;
    Number8[11][20] = 4'hF;
    Number8[12][20] = 4'hF;
    Number8[13][20] = 4'hF;
    Number8[14][20] = 4'hF;
    Number8[15][20] = 4'hD;
    Number8[16][20] = 4'hC;
    Number8[17][20] = 4'hC;
    Number8[18][20] = 4'hC;
    Number8[19][20] = 4'hC;
    Number8[20][20] = 4'hD;
    Number8[21][20] = 4'hF;
    Number8[22][20] = 4'hF;
    Number8[0][21] = 4'hF;
    Number8[1][21] = 4'hF;
    Number8[2][21] = 4'hE;
    Number8[3][21] = 4'hC;
    Number8[4][21] = 4'hC;
    Number8[5][21] = 4'hC;
    Number8[6][21] = 4'hC;
    Number8[7][21] = 4'hC;
    Number8[8][21] = 4'hE;
    Number8[9][21] = 4'hF;
    Number8[10][21] = 4'hF;
    Number8[11][21] = 4'hF;
    Number8[12][21] = 4'hF;
    Number8[13][21] = 4'hF;
    Number8[14][21] = 4'hF;
    Number8[15][21] = 4'hC;
    Number8[16][21] = 4'hC;
    Number8[17][21] = 4'hC;
    Number8[18][21] = 4'hC;
    Number8[19][21] = 4'hC;
    Number8[20][21] = 4'hD;
    Number8[21][21] = 4'hF;
    Number8[22][21] = 4'hF;
    Number8[0][22] = 4'hF;
    Number8[1][22] = 4'hF;
    Number8[2][22] = 4'hE;
    Number8[3][22] = 4'hC;
    Number8[4][22] = 4'hC;
    Number8[5][22] = 4'hC;
    Number8[6][22] = 4'hC;
    Number8[7][22] = 4'hC;
    Number8[8][22] = 4'hC;
    Number8[9][22] = 4'hD;
    Number8[10][22] = 4'hE;
    Number8[11][22] = 4'hF;
    Number8[12][22] = 4'hE;
    Number8[13][22] = 4'hD;
    Number8[14][22] = 4'hC;
    Number8[15][22] = 4'hC;
    Number8[16][22] = 4'hC;
    Number8[17][22] = 4'hC;
    Number8[18][22] = 4'hC;
    Number8[19][22] = 4'hC;
    Number8[20][22] = 4'hE;
    Number8[21][22] = 4'hF;
    Number8[22][22] = 4'hF;
    Number8[0][23] = 4'hF;
    Number8[1][23] = 4'hF;
    Number8[2][23] = 4'hF;
    Number8[3][23] = 4'hC;
    Number8[4][23] = 4'hC;
    Number8[5][23] = 4'hC;
    Number8[6][23] = 4'hC;
    Number8[7][23] = 4'hC;
    Number8[8][23] = 4'hC;
    Number8[9][23] = 4'hC;
    Number8[10][23] = 4'hC;
    Number8[11][23] = 4'hC;
    Number8[12][23] = 4'hC;
    Number8[13][23] = 4'hC;
    Number8[14][23] = 4'hC;
    Number8[15][23] = 4'hC;
    Number8[16][23] = 4'hC;
    Number8[17][23] = 4'hC;
    Number8[18][23] = 4'hC;
    Number8[19][23] = 4'hD;
    Number8[20][23] = 4'hF;
    Number8[21][23] = 4'hF;
    Number8[22][23] = 4'hF;
    Number8[0][24] = 4'hF;
    Number8[1][24] = 4'hF;
    Number8[2][24] = 4'hF;
    Number8[3][24] = 4'hE;
    Number8[4][24] = 4'hC;
    Number8[5][24] = 4'hC;
    Number8[6][24] = 4'hC;
    Number8[7][24] = 4'hC;
    Number8[8][24] = 4'hC;
    Number8[9][24] = 4'hC;
    Number8[10][24] = 4'hC;
    Number8[11][24] = 4'hC;
    Number8[12][24] = 4'hC;
    Number8[13][24] = 4'hC;
    Number8[14][24] = 4'hC;
    Number8[15][24] = 4'hC;
    Number8[16][24] = 4'hC;
    Number8[17][24] = 4'hC;
    Number8[18][24] = 4'hC;
    Number8[19][24] = 4'hE;
    Number8[20][24] = 4'hF;
    Number8[21][24] = 4'hF;
    Number8[22][24] = 4'hF;
    Number8[0][25] = 4'hF;
    Number8[1][25] = 4'hF;
    Number8[2][25] = 4'hF;
    Number8[3][25] = 4'hF;
    Number8[4][25] = 4'hE;
    Number8[5][25] = 4'hC;
    Number8[6][25] = 4'hC;
    Number8[7][25] = 4'hC;
    Number8[8][25] = 4'hC;
    Number8[9][25] = 4'hC;
    Number8[10][25] = 4'hC;
    Number8[11][25] = 4'hC;
    Number8[12][25] = 4'hC;
    Number8[13][25] = 4'hC;
    Number8[14][25] = 4'hC;
    Number8[15][25] = 4'hC;
    Number8[16][25] = 4'hC;
    Number8[17][25] = 4'hD;
    Number8[18][25] = 4'hE;
    Number8[19][25] = 4'hF;
    Number8[20][25] = 4'hF;
    Number8[21][25] = 4'hF;
    Number8[22][25] = 4'hF;
    Number8[0][26] = 4'hF;
    Number8[1][26] = 4'hF;
    Number8[2][26] = 4'hF;
    Number8[3][26] = 4'hF;
    Number8[4][26] = 4'hF;
    Number8[5][26] = 4'hF;
    Number8[6][26] = 4'hE;
    Number8[7][26] = 4'hD;
    Number8[8][26] = 4'hC;
    Number8[9][26] = 4'hC;
    Number8[10][26] = 4'hC;
    Number8[11][26] = 4'hC;
    Number8[12][26] = 4'hC;
    Number8[13][26] = 4'hC;
    Number8[14][26] = 4'hC;
    Number8[15][26] = 4'hD;
    Number8[16][26] = 4'hE;
    Number8[17][26] = 4'hF;
    Number8[18][26] = 4'hF;
    Number8[19][26] = 4'hF;
    Number8[20][26] = 4'hF;
    Number8[21][26] = 4'hF;
    Number8[22][26] = 4'hF;
    Number8[0][27] = 4'hF;
    Number8[1][27] = 4'hF;
    Number8[2][27] = 4'hF;
    Number8[3][27] = 4'hF;
    Number8[4][27] = 4'hF;
    Number8[5][27] = 4'hF;
    Number8[6][27] = 4'hF;
    Number8[7][27] = 4'hF;
    Number8[8][27] = 4'hF;
    Number8[9][27] = 4'hF;
    Number8[10][27] = 4'hF;
    Number8[11][27] = 4'hF;
    Number8[12][27] = 4'hF;
    Number8[13][27] = 4'hF;
    Number8[14][27] = 4'hF;
    Number8[15][27] = 4'hF;
    Number8[16][27] = 4'hF;
    Number8[17][27] = 4'hF;
    Number8[18][27] = 4'hF;
    Number8[19][27] = 4'hF;
    Number8[20][27] = 4'hF;
    Number8[21][27] = 4'hF;
    Number8[22][27] = 4'hF;
    Number8[0][28] = 4'hF;
    Number8[1][28] = 4'hF;
    Number8[2][28] = 4'hF;
    Number8[3][28] = 4'hF;
    Number8[4][28] = 4'hF;
    Number8[5][28] = 4'hF;
    Number8[6][28] = 4'hF;
    Number8[7][28] = 4'hF;
    Number8[8][28] = 4'hF;
    Number8[9][28] = 4'hF;
    Number8[10][28] = 4'hF;
    Number8[11][28] = 4'hF;
    Number8[12][28] = 4'hF;
    Number8[13][28] = 4'hF;
    Number8[14][28] = 4'hF;
    Number8[15][28] = 4'hF;
    Number8[16][28] = 4'hF;
    Number8[17][28] = 4'hF;
    Number8[18][28] = 4'hF;
    Number8[19][28] = 4'hF;
    Number8[20][28] = 4'hF;
    Number8[21][28] = 4'hF;
    Number8[22][28] = 4'hF;

// Number 9
    Number9[0][0] = 4'hF;
    Number9[1][0] = 4'hF;
    Number9[2][0] = 4'hF;
    Number9[3][0] = 4'hF;
    Number9[4][0] = 4'hF;
    Number9[5][0] = 4'hF;
    Number9[6][0] = 4'hF;
    Number9[7][0] = 4'hF;
    Number9[8][0] = 4'hF;
    Number9[9][0] = 4'hF;
    Number9[10][0] = 4'hF;
    Number9[11][0] = 4'hF;
    Number9[12][0] = 4'hF;
    Number9[13][0] = 4'hF;
    Number9[14][0] = 4'hF;
    Number9[15][0] = 4'hF;
    Number9[16][0] = 4'hF;
    Number9[17][0] = 4'hF;
    Number9[18][0] = 4'hF;
    Number9[19][0] = 4'hF;
    Number9[20][0] = 4'hF;
    Number9[21][0] = 4'hF;
    Number9[22][0] = 4'hF;
    Number9[0][1] = 4'hF;
    Number9[1][1] = 4'hF;
    Number9[2][1] = 4'hF;
    Number9[3][1] = 4'hF;
    Number9[4][1] = 4'hF;
    Number9[5][1] = 4'hF;
    Number9[6][1] = 4'hF;
    Number9[7][1] = 4'hF;
    Number9[8][1] = 4'hF;
    Number9[9][1] = 4'hF;
    Number9[10][1] = 4'hF;
    Number9[11][1] = 4'hF;
    Number9[12][1] = 4'hF;
    Number9[13][1] = 4'hF;
    Number9[14][1] = 4'hF;
    Number9[15][1] = 4'hF;
    Number9[16][1] = 4'hF;
    Number9[17][1] = 4'hF;
    Number9[18][1] = 4'hF;
    Number9[19][1] = 4'hF;
    Number9[20][1] = 4'hF;
    Number9[21][1] = 4'hF;
    Number9[22][1] = 4'hF;
    Number9[0][2] = 4'hF;
    Number9[1][2] = 4'hF;
    Number9[2][2] = 4'hF;
    Number9[3][2] = 4'hF;
    Number9[4][2] = 4'hF;
    Number9[5][2] = 4'hF;
    Number9[6][2] = 4'hF;
    Number9[7][2] = 4'hE;
    Number9[8][2] = 4'hD;
    Number9[9][2] = 4'hC;
    Number9[10][2] = 4'hC;
    Number9[11][2] = 4'hC;
    Number9[12][2] = 4'hC;
    Number9[13][2] = 4'hC;
    Number9[14][2] = 4'hD;
    Number9[15][2] = 4'hD;
    Number9[16][2] = 4'hF;
    Number9[17][2] = 4'hF;
    Number9[18][2] = 4'hF;
    Number9[19][2] = 4'hF;
    Number9[20][2] = 4'hF;
    Number9[21][2] = 4'hF;
    Number9[22][2] = 4'hF;
    Number9[0][3] = 4'hF;
    Number9[1][3] = 4'hF;
    Number9[2][3] = 4'hF;
    Number9[3][3] = 4'hF;
    Number9[4][3] = 4'hF;
    Number9[5][3] = 4'hE;
    Number9[6][3] = 4'hC;
    Number9[7][3] = 4'hC;
    Number9[8][3] = 4'hC;
    Number9[9][3] = 4'hC;
    Number9[10][3] = 4'hC;
    Number9[11][3] = 4'hC;
    Number9[12][3] = 4'hC;
    Number9[13][3] = 4'hC;
    Number9[14][3] = 4'hC;
    Number9[15][3] = 4'hC;
    Number9[16][3] = 4'hC;
    Number9[17][3] = 4'hE;
    Number9[18][3] = 4'hF;
    Number9[19][3] = 4'hF;
    Number9[20][3] = 4'hF;
    Number9[21][3] = 4'hF;
    Number9[22][3] = 4'hF;
    Number9[0][4] = 4'hF;
    Number9[1][4] = 4'hF;
    Number9[2][4] = 4'hF;
    Number9[3][4] = 4'hF;
    Number9[4][4] = 4'hE;
    Number9[5][4] = 4'hC;
    Number9[6][4] = 4'hC;
    Number9[7][4] = 4'hC;
    Number9[8][4] = 4'hC;
    Number9[9][4] = 4'hC;
    Number9[10][4] = 4'hC;
    Number9[11][4] = 4'hC;
    Number9[12][4] = 4'hC;
    Number9[13][4] = 4'hC;
    Number9[14][4] = 4'hC;
    Number9[15][4] = 4'hC;
    Number9[16][4] = 4'hC;
    Number9[17][4] = 4'hC;
    Number9[18][4] = 4'hE;
    Number9[19][4] = 4'hF;
    Number9[20][4] = 4'hF;
    Number9[21][4] = 4'hF;
    Number9[22][4] = 4'hF;
    Number9[0][5] = 4'hF;
    Number9[1][5] = 4'hF;
    Number9[2][5] = 4'hF;
    Number9[3][5] = 4'hF;
    Number9[4][5] = 4'hC;
    Number9[5][5] = 4'hC;
    Number9[6][5] = 4'hC;
    Number9[7][5] = 4'hC;
    Number9[8][5] = 4'hC;
    Number9[9][5] = 4'hC;
    Number9[10][5] = 4'hC;
    Number9[11][5] = 4'hC;
    Number9[12][5] = 4'hC;
    Number9[13][5] = 4'hC;
    Number9[14][5] = 4'hC;
    Number9[15][5] = 4'hC;
    Number9[16][5] = 4'hC;
    Number9[17][5] = 4'hC;
    Number9[18][5] = 4'hD;
    Number9[19][5] = 4'hF;
    Number9[20][5] = 4'hF;
    Number9[21][5] = 4'hF;
    Number9[22][5] = 4'hF;
    Number9[0][6] = 4'hF;
    Number9[1][6] = 4'hF;
    Number9[2][6] = 4'hF;
    Number9[3][6] = 4'hD;
    Number9[4][6] = 4'hC;
    Number9[5][6] = 4'hC;
    Number9[6][6] = 4'hC;
    Number9[7][6] = 4'hC;
    Number9[8][6] = 4'hC;
    Number9[9][6] = 4'hD;
    Number9[10][6] = 4'hE;
    Number9[11][6] = 4'hF;
    Number9[12][6] = 4'hE;
    Number9[13][6] = 4'hD;
    Number9[14][6] = 4'hC;
    Number9[15][6] = 4'hC;
    Number9[16][6] = 4'hC;
    Number9[17][6] = 4'hC;
    Number9[18][6] = 4'hC;
    Number9[19][6] = 4'hE;
    Number9[20][6] = 4'hF;
    Number9[21][6] = 4'hF;
    Number9[22][6] = 4'hF;
    Number9[0][7] = 4'hF;
    Number9[1][7] = 4'hF;
    Number9[2][7] = 4'hF;
    Number9[3][7] = 4'hC;
    Number9[4][7] = 4'hC;
    Number9[5][7] = 4'hC;
    Number9[6][7] = 4'hC;
    Number9[7][7] = 4'hC;
    Number9[8][7] = 4'hD;
    Number9[9][7] = 4'hF;
    Number9[10][7] = 4'hF;
    Number9[11][7] = 4'hF;
    Number9[12][7] = 4'hF;
    Number9[13][7] = 4'hF;
    Number9[14][7] = 4'hC;
    Number9[15][7] = 4'hC;
    Number9[16][7] = 4'hC;
    Number9[17][7] = 4'hC;
    Number9[18][7] = 4'hC;
    Number9[19][7] = 4'hD;
    Number9[20][7] = 4'hF;
    Number9[21][7] = 4'hF;
    Number9[22][7] = 4'hF;
    Number9[0][8] = 4'hF;
    Number9[1][8] = 4'hF;
    Number9[2][8] = 4'hF;
    Number9[3][8] = 4'hC;
    Number9[4][8] = 4'hC;
    Number9[5][8] = 4'hC;
    Number9[6][8] = 4'hC;
    Number9[7][8] = 4'hC;
    Number9[8][8] = 4'hE;
    Number9[9][8] = 4'hF;
    Number9[10][8] = 4'hF;
    Number9[11][8] = 4'hF;
    Number9[12][8] = 4'hF;
    Number9[13][8] = 4'hF;
    Number9[14][8] = 4'hD;
    Number9[15][8] = 4'hC;
    Number9[16][8] = 4'hC;
    Number9[17][8] = 4'hC;
    Number9[18][8] = 4'hC;
    Number9[19][8] = 4'hC;
    Number9[20][8] = 4'hF;
    Number9[21][8] = 4'hF;
    Number9[22][8] = 4'hF;
    Number9[0][9] = 4'hF;
    Number9[1][9] = 4'hF;
    Number9[2][9] = 4'hE;
    Number9[3][9] = 4'hC;
    Number9[4][9] = 4'hC;
    Number9[5][9] = 4'hC;
    Number9[6][9] = 4'hC;
    Number9[7][9] = 4'hC;
    Number9[8][9] = 4'hF;
    Number9[9][9] = 4'hF;
    Number9[10][9] = 4'hF;
    Number9[11][9] = 4'hF;
    Number9[12][9] = 4'hF;
    Number9[13][9] = 4'hF;
    Number9[14][9] = 4'hE;
    Number9[15][9] = 4'hC;
    Number9[16][9] = 4'hC;
    Number9[17][9] = 4'hC;
    Number9[18][9] = 4'hC;
    Number9[19][9] = 4'hC;
    Number9[20][9] = 4'hF;
    Number9[21][9] = 4'hF;
    Number9[22][9] = 4'hF;
    Number9[0][10] = 4'hF;
    Number9[1][10] = 4'hF;
    Number9[2][10] = 4'hE;
    Number9[3][10] = 4'hC;
    Number9[4][10] = 4'hC;
    Number9[5][10] = 4'hC;
    Number9[6][10] = 4'hC;
    Number9[7][10] = 4'hC;
    Number9[8][10] = 4'hF;
    Number9[9][10] = 4'hF;
    Number9[10][10] = 4'hF;
    Number9[11][10] = 4'hF;
    Number9[12][10] = 4'hF;
    Number9[13][10] = 4'hF;
    Number9[14][10] = 4'hF;
    Number9[15][10] = 4'hC;
    Number9[16][10] = 4'hC;
    Number9[17][10] = 4'hC;
    Number9[18][10] = 4'hC;
    Number9[19][10] = 4'hC;
    Number9[20][10] = 4'hE;
    Number9[21][10] = 4'hF;
    Number9[22][10] = 4'hF;
    Number9[0][11] = 4'hF;
    Number9[1][11] = 4'hF;
    Number9[2][11] = 4'hE;
    Number9[3][11] = 4'hC;
    Number9[4][11] = 4'hC;
    Number9[5][11] = 4'hC;
    Number9[6][11] = 4'hC;
    Number9[7][11] = 4'hC;
    Number9[8][11] = 4'hF;
    Number9[9][11] = 4'hF;
    Number9[10][11] = 4'hF;
    Number9[11][11] = 4'hF;
    Number9[12][11] = 4'hF;
    Number9[13][11] = 4'hF;
    Number9[14][11] = 4'hF;
    Number9[15][11] = 4'hC;
    Number9[16][11] = 4'hC;
    Number9[17][11] = 4'hC;
    Number9[18][11] = 4'hC;
    Number9[19][11] = 4'hC;
    Number9[20][11] = 4'hE;
    Number9[21][11] = 4'hF;
    Number9[22][11] = 4'hF;
    Number9[0][12] = 4'hF;
    Number9[1][12] = 4'hF;
    Number9[2][12] = 4'hF;
    Number9[3][12] = 4'hC;
    Number9[4][12] = 4'hC;
    Number9[5][12] = 4'hC;
    Number9[6][12] = 4'hC;
    Number9[7][12] = 4'hC;
    Number9[8][12] = 4'hD;
    Number9[9][12] = 4'hF;
    Number9[10][12] = 4'hF;
    Number9[11][12] = 4'hF;
    Number9[12][12] = 4'hF;
    Number9[13][12] = 4'hF;
    Number9[14][12] = 4'hF;
    Number9[15][12] = 4'hC;
    Number9[16][12] = 4'hC;
    Number9[17][12] = 4'hC;
    Number9[18][12] = 4'hC;
    Number9[19][12] = 4'hC;
    Number9[20][12] = 4'hE;
    Number9[21][12] = 4'hF;
    Number9[22][12] = 4'hF;
    Number9[0][13] = 4'hF;
    Number9[1][13] = 4'hF;
    Number9[2][13] = 4'hF;
    Number9[3][13] = 4'hC;
    Number9[4][13] = 4'hC;
    Number9[5][13] = 4'hC;
    Number9[6][13] = 4'hC;
    Number9[7][13] = 4'hC;
    Number9[8][13] = 4'hC;
    Number9[9][13] = 4'hD;
    Number9[10][13] = 4'hE;
    Number9[11][13] = 4'hF;
    Number9[12][13] = 4'hE;
    Number9[13][13] = 4'hD;
    Number9[14][13] = 4'hC;
    Number9[15][13] = 4'hC;
    Number9[16][13] = 4'hC;
    Number9[17][13] = 4'hC;
    Number9[18][13] = 4'hC;
    Number9[19][13] = 4'hC;
    Number9[20][13] = 4'hE;
    Number9[21][13] = 4'hF;
    Number9[22][13] = 4'hF;
    Number9[0][14] = 4'hF;
    Number9[1][14] = 4'hF;
    Number9[2][14] = 4'hF;
    Number9[3][14] = 4'hD;
    Number9[4][14] = 4'hC;
    Number9[5][14] = 4'hC;
    Number9[6][14] = 4'hC;
    Number9[7][14] = 4'hC;
    Number9[8][14] = 4'hC;
    Number9[9][14] = 4'hC;
    Number9[10][14] = 4'hC;
    Number9[11][14] = 4'hC;
    Number9[12][14] = 4'hC;
    Number9[13][14] = 4'hC;
    Number9[14][14] = 4'hC;
    Number9[15][14] = 4'hC;
    Number9[16][14] = 4'hC;
    Number9[17][14] = 4'hC;
    Number9[18][14] = 4'hC;
    Number9[19][14] = 4'hC;
    Number9[20][14] = 4'hE;
    Number9[21][14] = 4'hF;
    Number9[22][14] = 4'hF;
    Number9[0][15] = 4'hF;
    Number9[1][15] = 4'hF;
    Number9[2][15] = 4'hF;
    Number9[3][15] = 4'hF;
    Number9[4][15] = 4'hC;
    Number9[5][15] = 4'hC;
    Number9[6][15] = 4'hC;
    Number9[7][15] = 4'hC;
    Number9[8][15] = 4'hC;
    Number9[9][15] = 4'hC;
    Number9[10][15] = 4'hC;
    Number9[11][15] = 4'hC;
    Number9[12][15] = 4'hC;
    Number9[13][15] = 4'hC;
    Number9[14][15] = 4'hC;
    Number9[15][15] = 4'hC;
    Number9[16][15] = 4'hC;
    Number9[17][15] = 4'hC;
    Number9[18][15] = 4'hC;
    Number9[19][15] = 4'hC;
    Number9[20][15] = 4'hE;
    Number9[21][15] = 4'hF;
    Number9[22][15] = 4'hF;
    Number9[0][16] = 4'hF;
    Number9[1][16] = 4'hF;
    Number9[2][16] = 4'hF;
    Number9[3][16] = 4'hF;
    Number9[4][16] = 4'hE;
    Number9[5][16] = 4'hC;
    Number9[6][16] = 4'hC;
    Number9[7][16] = 4'hC;
    Number9[8][16] = 4'hC;
    Number9[9][16] = 4'hC;
    Number9[10][16] = 4'hC;
    Number9[11][16] = 4'hC;
    Number9[12][16] = 4'hC;
    Number9[13][16] = 4'hC;
    Number9[14][16] = 4'hC;
    Number9[15][16] = 4'hC;
    Number9[16][16] = 4'hC;
    Number9[17][16] = 4'hC;
    Number9[18][16] = 4'hC;
    Number9[19][16] = 4'hC;
    Number9[20][16] = 4'hE;
    Number9[21][16] = 4'hF;
    Number9[22][16] = 4'hF;
    Number9[0][17] = 4'hF;
    Number9[1][17] = 4'hF;
    Number9[2][17] = 4'hF;
    Number9[3][17] = 4'hF;
    Number9[4][17] = 4'hF;
    Number9[5][17] = 4'hF;
    Number9[6][17] = 4'hD;
    Number9[7][17] = 4'hD;
    Number9[8][17] = 4'hC;
    Number9[9][17] = 4'hC;
    Number9[10][17] = 4'hC;
    Number9[11][17] = 4'hC;
    Number9[12][17] = 4'hC;
    Number9[13][17] = 4'hD;
    Number9[14][17] = 4'hE;
    Number9[15][17] = 4'hC;
    Number9[16][17] = 4'hC;
    Number9[17][17] = 4'hC;
    Number9[18][17] = 4'hC;
    Number9[19][17] = 4'hC;
    Number9[20][17] = 4'hF;
    Number9[21][17] = 4'hF;
    Number9[22][17] = 4'hF;
    Number9[0][18] = 4'hF;
    Number9[1][18] = 4'hF;
    Number9[2][18] = 4'hF;
    Number9[3][18] = 4'hF;
    Number9[4][18] = 4'hF;
    Number9[5][18] = 4'hF;
    Number9[6][18] = 4'hF;
    Number9[7][18] = 4'hF;
    Number9[8][18] = 4'hF;
    Number9[9][18] = 4'hF;
    Number9[10][18] = 4'hF;
    Number9[11][18] = 4'hF;
    Number9[12][18] = 4'hF;
    Number9[13][18] = 4'hF;
    Number9[14][18] = 4'hF;
    Number9[15][18] = 4'hC;
    Number9[16][18] = 4'hC;
    Number9[17][18] = 4'hC;
    Number9[18][18] = 4'hC;
    Number9[19][18] = 4'hC;
    Number9[20][18] = 4'hF;
    Number9[21][18] = 4'hF;
    Number9[22][18] = 4'hF;
    Number9[0][19] = 4'hF;
    Number9[1][19] = 4'hF;
    Number9[2][19] = 4'hF;
    Number9[3][19] = 4'hF;
    Number9[4][19] = 4'hF;
    Number9[5][19] = 4'hF;
    Number9[6][19] = 4'hF;
    Number9[7][19] = 4'hF;
    Number9[8][19] = 4'hF;
    Number9[9][19] = 4'hF;
    Number9[10][19] = 4'hF;
    Number9[11][19] = 4'hF;
    Number9[12][19] = 4'hF;
    Number9[13][19] = 4'hF;
    Number9[14][19] = 4'hD;
    Number9[15][19] = 4'hC;
    Number9[16][19] = 4'hC;
    Number9[17][19] = 4'hC;
    Number9[18][19] = 4'hC;
    Number9[19][19] = 4'hD;
    Number9[20][19] = 4'hF;
    Number9[21][19] = 4'hF;
    Number9[22][19] = 4'hF;
    Number9[0][20] = 4'hF;
    Number9[1][20] = 4'hF;
    Number9[2][20] = 4'hF;
    Number9[3][20] = 4'hF;
    Number9[4][20] = 4'hF;
    Number9[5][20] = 4'hF;
    Number9[6][20] = 4'hF;
    Number9[7][20] = 4'hF;
    Number9[8][20] = 4'hF;
    Number9[9][20] = 4'hF;
    Number9[10][20] = 4'hF;
    Number9[11][20] = 4'hF;
    Number9[12][20] = 4'hF;
    Number9[13][20] = 4'hF;
    Number9[14][20] = 4'hC;
    Number9[15][20] = 4'hC;
    Number9[16][20] = 4'hC;
    Number9[17][20] = 4'hC;
    Number9[18][20] = 4'hC;
    Number9[19][20] = 4'hE;
    Number9[20][20] = 4'hF;
    Number9[21][20] = 4'hF;
    Number9[22][20] = 4'hF;
    Number9[0][21] = 4'hF;
    Number9[1][21] = 4'hF;
    Number9[2][21] = 4'hF;
    Number9[3][21] = 4'hF;
    Number9[4][21] = 4'hF;
    Number9[5][21] = 4'hF;
    Number9[6][21] = 4'hF;
    Number9[7][21] = 4'hF;
    Number9[8][21] = 4'hF;
    Number9[9][21] = 4'hF;
    Number9[10][21] = 4'hF;
    Number9[11][21] = 4'hF;
    Number9[12][21] = 4'hF;
    Number9[13][21] = 4'hD;
    Number9[14][21] = 4'hC;
    Number9[15][21] = 4'hC;
    Number9[16][21] = 4'hC;
    Number9[17][21] = 4'hC;
    Number9[18][21] = 4'hC;
    Number9[19][21] = 4'hF;
    Number9[20][21] = 4'hF;
    Number9[21][21] = 4'hF;
    Number9[22][21] = 4'hF;
    Number9[0][22] = 4'hF;
    Number9[1][22] = 4'hF;
    Number9[2][22] = 4'hF;
    Number9[3][22] = 4'hE;
    Number9[4][22] = 4'hC;
    Number9[5][22] = 4'hD;
    Number9[6][22] = 4'hD;
    Number9[7][22] = 4'hE;
    Number9[8][22] = 4'hE;
    Number9[9][22] = 4'hF;
    Number9[10][22] = 4'hE;
    Number9[11][22] = 4'hD;
    Number9[12][22] = 4'hC;
    Number9[13][22] = 4'hC;
    Number9[14][22] = 4'hC;
    Number9[15][22] = 4'hC;
    Number9[16][22] = 4'hC;
    Number9[17][22] = 4'hC;
    Number9[18][22] = 4'hE;
    Number9[19][22] = 4'hF;
    Number9[20][22] = 4'hF;
    Number9[21][22] = 4'hF;
    Number9[22][22] = 4'hF;
    Number9[0][23] = 4'hF;
    Number9[1][23] = 4'hF;
    Number9[2][23] = 4'hF;
    Number9[3][23] = 4'hD;
    Number9[4][23] = 4'hC;
    Number9[5][23] = 4'hC;
    Number9[6][23] = 4'hC;
    Number9[7][23] = 4'hC;
    Number9[8][23] = 4'hC;
    Number9[9][23] = 4'hC;
    Number9[10][23] = 4'hC;
    Number9[11][23] = 4'hC;
    Number9[12][23] = 4'hC;
    Number9[13][23] = 4'hC;
    Number9[14][23] = 4'hC;
    Number9[15][23] = 4'hC;
    Number9[16][23] = 4'hC;
    Number9[17][23] = 4'hD;
    Number9[18][23] = 4'hF;
    Number9[19][23] = 4'hF;
    Number9[20][23] = 4'hF;
    Number9[21][23] = 4'hF;
    Number9[22][23] = 4'hF;
    Number9[0][24] = 4'hF;
    Number9[1][24] = 4'hF;
    Number9[2][24] = 4'hF;
    Number9[3][24] = 4'hE;
    Number9[4][24] = 4'hC;
    Number9[5][24] = 4'hC;
    Number9[6][24] = 4'hC;
    Number9[7][24] = 4'hC;
    Number9[8][24] = 4'hC;
    Number9[9][24] = 4'hC;
    Number9[10][24] = 4'hC;
    Number9[11][24] = 4'hC;
    Number9[12][24] = 4'hC;
    Number9[13][24] = 4'hC;
    Number9[14][24] = 4'hC;
    Number9[15][24] = 4'hC;
    Number9[16][24] = 4'hD;
    Number9[17][24] = 4'hF;
    Number9[18][24] = 4'hF;
    Number9[19][24] = 4'hF;
    Number9[20][24] = 4'hF;
    Number9[21][24] = 4'hF;
    Number9[22][24] = 4'hF;
    Number9[0][25] = 4'hF;
    Number9[1][25] = 4'hF;
    Number9[2][25] = 4'hF;
    Number9[3][25] = 4'hE;
    Number9[4][25] = 4'hC;
    Number9[5][25] = 4'hC;
    Number9[6][25] = 4'hC;
    Number9[7][25] = 4'hC;
    Number9[8][25] = 4'hC;
    Number9[9][25] = 4'hC;
    Number9[10][25] = 4'hC;
    Number9[11][25] = 4'hC;
    Number9[12][25] = 4'hC;
    Number9[13][25] = 4'hC;
    Number9[14][25] = 4'hC;
    Number9[15][25] = 4'hD;
    Number9[16][25] = 4'hF;
    Number9[17][25] = 4'hF;
    Number9[18][25] = 4'hF;
    Number9[19][25] = 4'hF;
    Number9[20][25] = 4'hF;
    Number9[21][25] = 4'hF;
    Number9[22][25] = 4'hF;
    Number9[0][26] = 4'hF;
    Number9[1][26] = 4'hF;
    Number9[2][26] = 4'hF;
    Number9[3][26] = 4'hF;
    Number9[4][26] = 4'hE;
    Number9[5][26] = 4'hD;
    Number9[6][26] = 4'hD;
    Number9[7][26] = 4'hC;
    Number9[8][26] = 4'hC;
    Number9[9][26] = 4'hC;
    Number9[10][26] = 4'hC;
    Number9[11][26] = 4'hC;
    Number9[12][26] = 4'hD;
    Number9[13][26] = 4'hD;
    Number9[14][26] = 4'hF;
    Number9[15][26] = 4'hF;
    Number9[16][26] = 4'hF;
    Number9[17][26] = 4'hF;
    Number9[18][26] = 4'hF;
    Number9[19][26] = 4'hF;
    Number9[20][26] = 4'hF;
    Number9[21][26] = 4'hF;
    Number9[22][26] = 4'hF;
    Number9[0][27] = 4'hF;
    Number9[1][27] = 4'hF;
    Number9[2][27] = 4'hF;
    Number9[3][27] = 4'hF;
    Number9[4][27] = 4'hF;
    Number9[5][27] = 4'hF;
    Number9[6][27] = 4'hF;
    Number9[7][27] = 4'hF;
    Number9[8][27] = 4'hF;
    Number9[9][27] = 4'hF;
    Number9[10][27] = 4'hF;
    Number9[11][27] = 4'hF;
    Number9[12][27] = 4'hF;
    Number9[13][27] = 4'hF;
    Number9[14][27] = 4'hF;
    Number9[15][27] = 4'hF;
    Number9[16][27] = 4'hF;
    Number9[17][27] = 4'hF;
    Number9[18][27] = 4'hF;
    Number9[19][27] = 4'hF;
    Number9[20][27] = 4'hF;
    Number9[21][27] = 4'hF;
    Number9[22][27] = 4'hF;
    Number9[0][28] = 4'hF;
    Number9[1][28] = 4'hF;
    Number9[2][28] = 4'hF;
    Number9[3][28] = 4'hF;
    Number9[4][28] = 4'hF;
    Number9[5][28] = 4'hF;
    Number9[6][28] = 4'hF;
    Number9[7][28] = 4'hF;
    Number9[8][28] = 4'hF;
    Number9[9][28] = 4'hF;
    Number9[10][28] = 4'hF;
    Number9[11][28] = 4'hF;
    Number9[12][28] = 4'hF;
    Number9[13][28] = 4'hF;
    Number9[14][28] = 4'hF;
    Number9[15][28] = 4'hF;
    Number9[16][28] = 4'hF;
    Number9[17][28] = 4'hF;
    Number9[18][28] = 4'hF;
    Number9[19][28] = 4'hF;
    Number9[20][28] = 4'hF;
    Number9[21][28] = 4'hF;
    Number9[22][28] = 4'hF;

end

endmodule
