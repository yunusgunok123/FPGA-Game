module Spaceship_init (
		output reg [3:0] SS0[0:47][0:47],
		output reg [3:0] SS1[0:47][0:47],
		output reg [3:0] SS2[0:47][0:47],
		output reg [3:0] SS3[0:47][0:47],
		output reg [3:0] SS4[0:47][0:47],
		output reg [3:0] SS5[0:47][0:47],
		output reg [3:0] SS6[0:47][0:47],
		output reg [3:0] SS7[0:47][0:47],
		output reg [3:0] SS8[0:47][0:47],
		output reg [3:0] SS9[0:47][0:47],
		output reg [3:0] SS10[0:47][0:47],
		output reg [3:0] SS11[0:47][0:47],
		output reg [3:0] SS12[0:47][0:47],
		output reg [3:0] SS13[0:47][0:47],
		output reg [3:0] SS14[0:47][0:47],
		output reg [3:0] SS15[0:47][0:47]
);
// Storing the pixel color information of Pictures of spaceships for each direction
initial begin

//SS 0
    SS0[0][0] = 4'h0;
    SS0[1][0] = 4'h0;
    SS0[2][0] = 4'h0;
    SS0[3][0] = 4'h0;
    SS0[4][0] = 4'h0;
    SS0[5][0] = 4'h0;
    SS0[6][0] = 4'h0;
    SS0[7][0] = 4'h0;
    SS0[8][0] = 4'h0;
    SS0[9][0] = 4'hD;
    SS0[10][0] = 4'hD;
    SS0[11][0] = 4'hD;
    SS0[12][0] = 4'h0;
    SS0[13][0] = 4'h0;
    SS0[14][0] = 4'h0;
    SS0[15][0] = 4'h0;
    SS0[16][0] = 4'h0;
    SS0[17][0] = 4'h0;
    SS0[18][0] = 4'h0;
    SS0[19][0] = 4'h0;
    SS0[20][0] = 4'h0;
    SS0[21][0] = 4'h0;
    SS0[22][0] = 4'h0;
    SS0[23][0] = 4'h0;
    SS0[24][0] = 4'h0;
    SS0[25][0] = 4'h0;
    SS0[26][0] = 4'h0;
    SS0[27][0] = 4'h0;
    SS0[28][0] = 4'h0;
    SS0[29][0] = 4'h0;
    SS0[30][0] = 4'h0;
    SS0[31][0] = 4'h0;
    SS0[32][0] = 4'h0;
    SS0[33][0] = 4'h0;
    SS0[34][0] = 4'h0;
    SS0[35][0] = 4'h0;
    SS0[36][0] = 4'hD;
    SS0[37][0] = 4'hD;
    SS0[38][0] = 4'hD;
    SS0[39][0] = 4'h0;
    SS0[40][0] = 4'h0;
    SS0[41][0] = 4'h0;
    SS0[42][0] = 4'h0;
    SS0[43][0] = 4'h0;
    SS0[44][0] = 4'h0;
    SS0[45][0] = 4'h0;
    SS0[46][0] = 4'h0;
    SS0[47][0] = 4'h0;
    SS0[0][1] = 4'h0;
    SS0[1][1] = 4'h0;
    SS0[2][1] = 4'h0;
    SS0[3][1] = 4'h0;
    SS0[4][1] = 4'h0;
    SS0[5][1] = 4'h0;
    SS0[6][1] = 4'h0;
    SS0[7][1] = 4'h0;
    SS0[8][1] = 4'h0;
    SS0[9][1] = 4'hD;
    SS0[10][1] = 4'hD;
    SS0[11][1] = 4'hD;
    SS0[12][1] = 4'h0;
    SS0[13][1] = 4'h0;
    SS0[14][1] = 4'h0;
    SS0[15][1] = 4'h0;
    SS0[16][1] = 4'h0;
    SS0[17][1] = 4'h0;
    SS0[18][1] = 4'h0;
    SS0[19][1] = 4'h0;
    SS0[20][1] = 4'h0;
    SS0[21][1] = 4'h0;
    SS0[22][1] = 4'h0;
    SS0[23][1] = 4'h0;
    SS0[24][1] = 4'h0;
    SS0[25][1] = 4'h0;
    SS0[26][1] = 4'h0;
    SS0[27][1] = 4'h0;
    SS0[28][1] = 4'h0;
    SS0[29][1] = 4'h0;
    SS0[30][1] = 4'h0;
    SS0[31][1] = 4'h0;
    SS0[32][1] = 4'h0;
    SS0[33][1] = 4'h0;
    SS0[34][1] = 4'h0;
    SS0[35][1] = 4'h0;
    SS0[36][1] = 4'hD;
    SS0[37][1] = 4'hD;
    SS0[38][1] = 4'hD;
    SS0[39][1] = 4'h0;
    SS0[40][1] = 4'h0;
    SS0[41][1] = 4'h0;
    SS0[42][1] = 4'h0;
    SS0[43][1] = 4'h0;
    SS0[44][1] = 4'h0;
    SS0[45][1] = 4'h0;
    SS0[46][1] = 4'h0;
    SS0[47][1] = 4'h0;
    SS0[0][2] = 4'h0;
    SS0[1][2] = 4'h0;
    SS0[2][2] = 4'h0;
    SS0[3][2] = 4'h0;
    SS0[4][2] = 4'h0;
    SS0[5][2] = 4'h0;
    SS0[6][2] = 4'h0;
    SS0[7][2] = 4'h0;
    SS0[8][2] = 4'h0;
    SS0[9][2] = 4'hD;
    SS0[10][2] = 4'hD;
    SS0[11][2] = 4'hD;
    SS0[12][2] = 4'h0;
    SS0[13][2] = 4'h0;
    SS0[14][2] = 4'h0;
    SS0[15][2] = 4'h0;
    SS0[16][2] = 4'h0;
    SS0[17][2] = 4'h0;
    SS0[18][2] = 4'h0;
    SS0[19][2] = 4'h0;
    SS0[20][2] = 4'h0;
    SS0[21][2] = 4'h0;
    SS0[22][2] = 4'h0;
    SS0[23][2] = 4'h0;
    SS0[24][2] = 4'h0;
    SS0[25][2] = 4'h0;
    SS0[26][2] = 4'h0;
    SS0[27][2] = 4'h0;
    SS0[28][2] = 4'h0;
    SS0[29][2] = 4'h0;
    SS0[30][2] = 4'h0;
    SS0[31][2] = 4'h0;
    SS0[32][2] = 4'h0;
    SS0[33][2] = 4'h0;
    SS0[34][2] = 4'h0;
    SS0[35][2] = 4'h0;
    SS0[36][2] = 4'hD;
    SS0[37][2] = 4'hD;
    SS0[38][2] = 4'hD;
    SS0[39][2] = 4'h0;
    SS0[40][2] = 4'h0;
    SS0[41][2] = 4'h0;
    SS0[42][2] = 4'h0;
    SS0[43][2] = 4'h0;
    SS0[44][2] = 4'h0;
    SS0[45][2] = 4'h0;
    SS0[46][2] = 4'h0;
    SS0[47][2] = 4'h0;
    SS0[0][3] = 4'h0;
    SS0[1][3] = 4'h0;
    SS0[2][3] = 4'h0;
    SS0[3][3] = 4'h0;
    SS0[4][3] = 4'h0;
    SS0[5][3] = 4'h0;
    SS0[6][3] = 4'h0;
    SS0[7][3] = 4'h0;
    SS0[8][3] = 4'h0;
    SS0[9][3] = 4'hC;
    SS0[10][3] = 4'hC;
    SS0[11][3] = 4'hC;
    SS0[12][3] = 4'hD;
    SS0[13][3] = 4'hD;
    SS0[14][3] = 4'hD;
    SS0[15][3] = 4'h0;
    SS0[16][3] = 4'h0;
    SS0[17][3] = 4'h0;
    SS0[18][3] = 4'h0;
    SS0[19][3] = 4'h0;
    SS0[20][3] = 4'h0;
    SS0[21][3] = 4'h0;
    SS0[22][3] = 4'h0;
    SS0[23][3] = 4'h0;
    SS0[24][3] = 4'h0;
    SS0[25][3] = 4'h0;
    SS0[26][3] = 4'h0;
    SS0[27][3] = 4'h0;
    SS0[28][3] = 4'h0;
    SS0[29][3] = 4'h0;
    SS0[30][3] = 4'h0;
    SS0[31][3] = 4'h0;
    SS0[32][3] = 4'h0;
    SS0[33][3] = 4'hD;
    SS0[34][3] = 4'hD;
    SS0[35][3] = 4'hD;
    SS0[36][3] = 4'hC;
    SS0[37][3] = 4'hC;
    SS0[38][3] = 4'hC;
    SS0[39][3] = 4'h0;
    SS0[40][3] = 4'h0;
    SS0[41][3] = 4'h0;
    SS0[42][3] = 4'h0;
    SS0[43][3] = 4'h0;
    SS0[44][3] = 4'h0;
    SS0[45][3] = 4'h0;
    SS0[46][3] = 4'h0;
    SS0[47][3] = 4'h0;
    SS0[0][4] = 4'h0;
    SS0[1][4] = 4'h0;
    SS0[2][4] = 4'h0;
    SS0[3][4] = 4'h0;
    SS0[4][4] = 4'h0;
    SS0[5][4] = 4'h0;
    SS0[6][4] = 4'h0;
    SS0[7][4] = 4'h0;
    SS0[8][4] = 4'h0;
    SS0[9][4] = 4'hC;
    SS0[10][4] = 4'hC;
    SS0[11][4] = 4'hC;
    SS0[12][4] = 4'hD;
    SS0[13][4] = 4'hD;
    SS0[14][4] = 4'hD;
    SS0[15][4] = 4'h0;
    SS0[16][4] = 4'h0;
    SS0[17][4] = 4'h0;
    SS0[18][4] = 4'h0;
    SS0[19][4] = 4'h0;
    SS0[20][4] = 4'h0;
    SS0[21][4] = 4'h0;
    SS0[22][4] = 4'h0;
    SS0[23][4] = 4'h0;
    SS0[24][4] = 4'h0;
    SS0[25][4] = 4'h0;
    SS0[26][4] = 4'h0;
    SS0[27][4] = 4'h0;
    SS0[28][4] = 4'h0;
    SS0[29][4] = 4'h0;
    SS0[30][4] = 4'h0;
    SS0[31][4] = 4'h0;
    SS0[32][4] = 4'h0;
    SS0[33][4] = 4'hD;
    SS0[34][4] = 4'hD;
    SS0[35][4] = 4'hD;
    SS0[36][4] = 4'hC;
    SS0[37][4] = 4'hC;
    SS0[38][4] = 4'hC;
    SS0[39][4] = 4'h0;
    SS0[40][4] = 4'h0;
    SS0[41][4] = 4'h0;
    SS0[42][4] = 4'h0;
    SS0[43][4] = 4'h0;
    SS0[44][4] = 4'h0;
    SS0[45][4] = 4'h0;
    SS0[46][4] = 4'h0;
    SS0[47][4] = 4'h0;
    SS0[0][5] = 4'h0;
    SS0[1][5] = 4'h0;
    SS0[2][5] = 4'h0;
    SS0[3][5] = 4'h0;
    SS0[4][5] = 4'h0;
    SS0[5][5] = 4'h0;
    SS0[6][5] = 4'h0;
    SS0[7][5] = 4'h0;
    SS0[8][5] = 4'h0;
    SS0[9][5] = 4'hC;
    SS0[10][5] = 4'hC;
    SS0[11][5] = 4'hC;
    SS0[12][5] = 4'hD;
    SS0[13][5] = 4'hD;
    SS0[14][5] = 4'hD;
    SS0[15][5] = 4'h0;
    SS0[16][5] = 4'h0;
    SS0[17][5] = 4'h0;
    SS0[18][5] = 4'h0;
    SS0[19][5] = 4'h0;
    SS0[20][5] = 4'h0;
    SS0[21][5] = 4'h0;
    SS0[22][5] = 4'h0;
    SS0[23][5] = 4'h0;
    SS0[24][5] = 4'h0;
    SS0[25][5] = 4'h0;
    SS0[26][5] = 4'h0;
    SS0[27][5] = 4'h0;
    SS0[28][5] = 4'h0;
    SS0[29][5] = 4'h0;
    SS0[30][5] = 4'h0;
    SS0[31][5] = 4'h0;
    SS0[32][5] = 4'h0;
    SS0[33][5] = 4'hD;
    SS0[34][5] = 4'hD;
    SS0[35][5] = 4'hD;
    SS0[36][5] = 4'hC;
    SS0[37][5] = 4'hC;
    SS0[38][5] = 4'hC;
    SS0[39][5] = 4'h0;
    SS0[40][5] = 4'h0;
    SS0[41][5] = 4'h0;
    SS0[42][5] = 4'h0;
    SS0[43][5] = 4'h0;
    SS0[44][5] = 4'h0;
    SS0[45][5] = 4'h0;
    SS0[46][5] = 4'h0;
    SS0[47][5] = 4'h0;
    SS0[0][6] = 4'h0;
    SS0[1][6] = 4'h0;
    SS0[2][6] = 4'h0;
    SS0[3][6] = 4'h0;
    SS0[4][6] = 4'h0;
    SS0[5][6] = 4'h0;
    SS0[6][6] = 4'h0;
    SS0[7][6] = 4'h0;
    SS0[8][6] = 4'h0;
    SS0[9][6] = 4'hC;
    SS0[10][6] = 4'hC;
    SS0[11][6] = 4'hC;
    SS0[12][6] = 4'hC;
    SS0[13][6] = 4'hC;
    SS0[14][6] = 4'hC;
    SS0[15][6] = 4'hE;
    SS0[16][6] = 4'hE;
    SS0[17][6] = 4'hE;
    SS0[18][6] = 4'h0;
    SS0[19][6] = 4'h0;
    SS0[20][6] = 4'h0;
    SS0[21][6] = 4'h0;
    SS0[22][6] = 4'h0;
    SS0[23][6] = 4'h0;
    SS0[24][6] = 4'h0;
    SS0[25][6] = 4'h0;
    SS0[26][6] = 4'h0;
    SS0[27][6] = 4'h0;
    SS0[28][6] = 4'h0;
    SS0[29][6] = 4'h0;
    SS0[30][6] = 4'hE;
    SS0[31][6] = 4'hE;
    SS0[32][6] = 4'hE;
    SS0[33][6] = 4'hC;
    SS0[34][6] = 4'hC;
    SS0[35][6] = 4'hC;
    SS0[36][6] = 4'hC;
    SS0[37][6] = 4'hC;
    SS0[38][6] = 4'hC;
    SS0[39][6] = 4'h0;
    SS0[40][6] = 4'h0;
    SS0[41][6] = 4'h0;
    SS0[42][6] = 4'h0;
    SS0[43][6] = 4'h0;
    SS0[44][6] = 4'h0;
    SS0[45][6] = 4'h0;
    SS0[46][6] = 4'h0;
    SS0[47][6] = 4'h0;
    SS0[0][7] = 4'h0;
    SS0[1][7] = 4'h0;
    SS0[2][7] = 4'h0;
    SS0[3][7] = 4'h0;
    SS0[4][7] = 4'h0;
    SS0[5][7] = 4'h0;
    SS0[6][7] = 4'h0;
    SS0[7][7] = 4'h0;
    SS0[8][7] = 4'h0;
    SS0[9][7] = 4'hC;
    SS0[10][7] = 4'hC;
    SS0[11][7] = 4'hC;
    SS0[12][7] = 4'hC;
    SS0[13][7] = 4'hC;
    SS0[14][7] = 4'hC;
    SS0[15][7] = 4'hE;
    SS0[16][7] = 4'hE;
    SS0[17][7] = 4'hE;
    SS0[18][7] = 4'h0;
    SS0[19][7] = 4'h0;
    SS0[20][7] = 4'h0;
    SS0[21][7] = 4'h0;
    SS0[22][7] = 4'h0;
    SS0[23][7] = 4'h0;
    SS0[24][7] = 4'h0;
    SS0[25][7] = 4'h0;
    SS0[26][7] = 4'h0;
    SS0[27][7] = 4'h0;
    SS0[28][7] = 4'h0;
    SS0[29][7] = 4'h0;
    SS0[30][7] = 4'hE;
    SS0[31][7] = 4'hE;
    SS0[32][7] = 4'hE;
    SS0[33][7] = 4'hC;
    SS0[34][7] = 4'hC;
    SS0[35][7] = 4'hC;
    SS0[36][7] = 4'hC;
    SS0[37][7] = 4'hC;
    SS0[38][7] = 4'hC;
    SS0[39][7] = 4'h0;
    SS0[40][7] = 4'h0;
    SS0[41][7] = 4'h0;
    SS0[42][7] = 4'h0;
    SS0[43][7] = 4'h0;
    SS0[44][7] = 4'h0;
    SS0[45][7] = 4'h0;
    SS0[46][7] = 4'h0;
    SS0[47][7] = 4'h0;
    SS0[0][8] = 4'h0;
    SS0[1][8] = 4'h0;
    SS0[2][8] = 4'h0;
    SS0[3][8] = 4'h0;
    SS0[4][8] = 4'h0;
    SS0[5][8] = 4'h0;
    SS0[6][8] = 4'h0;
    SS0[7][8] = 4'h0;
    SS0[8][8] = 4'h0;
    SS0[9][8] = 4'hC;
    SS0[10][8] = 4'hC;
    SS0[11][8] = 4'hC;
    SS0[12][8] = 4'hC;
    SS0[13][8] = 4'hC;
    SS0[14][8] = 4'hC;
    SS0[15][8] = 4'hE;
    SS0[16][8] = 4'hE;
    SS0[17][8] = 4'hE;
    SS0[18][8] = 4'h0;
    SS0[19][8] = 4'h0;
    SS0[20][8] = 4'h0;
    SS0[21][8] = 4'h0;
    SS0[22][8] = 4'h0;
    SS0[23][8] = 4'h0;
    SS0[24][8] = 4'h0;
    SS0[25][8] = 4'h0;
    SS0[26][8] = 4'h0;
    SS0[27][8] = 4'h0;
    SS0[28][8] = 4'h0;
    SS0[29][8] = 4'h0;
    SS0[30][8] = 4'hE;
    SS0[31][8] = 4'hE;
    SS0[32][8] = 4'hE;
    SS0[33][8] = 4'hC;
    SS0[34][8] = 4'hC;
    SS0[35][8] = 4'hC;
    SS0[36][8] = 4'hC;
    SS0[37][8] = 4'hC;
    SS0[38][8] = 4'hC;
    SS0[39][8] = 4'h0;
    SS0[40][8] = 4'h0;
    SS0[41][8] = 4'h0;
    SS0[42][8] = 4'h0;
    SS0[43][8] = 4'h0;
    SS0[44][8] = 4'h0;
    SS0[45][8] = 4'h0;
    SS0[46][8] = 4'h0;
    SS0[47][8] = 4'h0;
    SS0[0][9] = 4'h0;
    SS0[1][9] = 4'h0;
    SS0[2][9] = 4'h0;
    SS0[3][9] = 4'h0;
    SS0[4][9] = 4'h0;
    SS0[5][9] = 4'h0;
    SS0[6][9] = 4'h0;
    SS0[7][9] = 4'h0;
    SS0[8][9] = 4'h0;
    SS0[9][9] = 4'h0;
    SS0[10][9] = 4'h0;
    SS0[11][9] = 4'h0;
    SS0[12][9] = 4'hC;
    SS0[13][9] = 4'hC;
    SS0[14][9] = 4'hC;
    SS0[15][9] = 4'hD;
    SS0[16][9] = 4'hD;
    SS0[17][9] = 4'hD;
    SS0[18][9] = 4'hE;
    SS0[19][9] = 4'hE;
    SS0[20][9] = 4'hE;
    SS0[21][9] = 4'h0;
    SS0[22][9] = 4'h0;
    SS0[23][9] = 4'h0;
    SS0[24][9] = 4'h0;
    SS0[25][9] = 4'h0;
    SS0[26][9] = 4'h0;
    SS0[27][9] = 4'hE;
    SS0[28][9] = 4'hE;
    SS0[29][9] = 4'hE;
    SS0[30][9] = 4'hD;
    SS0[31][9] = 4'hD;
    SS0[32][9] = 4'hD;
    SS0[33][9] = 4'hC;
    SS0[34][9] = 4'hC;
    SS0[35][9] = 4'hC;
    SS0[36][9] = 4'h0;
    SS0[37][9] = 4'h0;
    SS0[38][9] = 4'h0;
    SS0[39][9] = 4'h0;
    SS0[40][9] = 4'h0;
    SS0[41][9] = 4'h0;
    SS0[42][9] = 4'h0;
    SS0[43][9] = 4'h0;
    SS0[44][9] = 4'h0;
    SS0[45][9] = 4'h0;
    SS0[46][9] = 4'h0;
    SS0[47][9] = 4'h0;
    SS0[0][10] = 4'h0;
    SS0[1][10] = 4'h0;
    SS0[2][10] = 4'h0;
    SS0[3][10] = 4'h0;
    SS0[4][10] = 4'h0;
    SS0[5][10] = 4'h0;
    SS0[6][10] = 4'h0;
    SS0[7][10] = 4'h0;
    SS0[8][10] = 4'h0;
    SS0[9][10] = 4'h0;
    SS0[10][10] = 4'h0;
    SS0[11][10] = 4'h0;
    SS0[12][10] = 4'hC;
    SS0[13][10] = 4'hC;
    SS0[14][10] = 4'hC;
    SS0[15][10] = 4'hD;
    SS0[16][10] = 4'hD;
    SS0[17][10] = 4'hD;
    SS0[18][10] = 4'hE;
    SS0[19][10] = 4'hE;
    SS0[20][10] = 4'hE;
    SS0[21][10] = 4'h0;
    SS0[22][10] = 4'h0;
    SS0[23][10] = 4'h0;
    SS0[24][10] = 4'h0;
    SS0[25][10] = 4'h0;
    SS0[26][10] = 4'h0;
    SS0[27][10] = 4'hE;
    SS0[28][10] = 4'hE;
    SS0[29][10] = 4'hE;
    SS0[30][10] = 4'hD;
    SS0[31][10] = 4'hD;
    SS0[32][10] = 4'hD;
    SS0[33][10] = 4'hC;
    SS0[34][10] = 4'hC;
    SS0[35][10] = 4'hC;
    SS0[36][10] = 4'h0;
    SS0[37][10] = 4'h0;
    SS0[38][10] = 4'h0;
    SS0[39][10] = 4'h0;
    SS0[40][10] = 4'h0;
    SS0[41][10] = 4'h0;
    SS0[42][10] = 4'h0;
    SS0[43][10] = 4'h0;
    SS0[44][10] = 4'h0;
    SS0[45][10] = 4'h0;
    SS0[46][10] = 4'h0;
    SS0[47][10] = 4'h0;
    SS0[0][11] = 4'h0;
    SS0[1][11] = 4'h0;
    SS0[2][11] = 4'h0;
    SS0[3][11] = 4'h0;
    SS0[4][11] = 4'h0;
    SS0[5][11] = 4'h0;
    SS0[6][11] = 4'h0;
    SS0[7][11] = 4'h0;
    SS0[8][11] = 4'h0;
    SS0[9][11] = 4'h0;
    SS0[10][11] = 4'h0;
    SS0[11][11] = 4'h0;
    SS0[12][11] = 4'hC;
    SS0[13][11] = 4'hC;
    SS0[14][11] = 4'hC;
    SS0[15][11] = 4'hD;
    SS0[16][11] = 4'hD;
    SS0[17][11] = 4'hD;
    SS0[18][11] = 4'hE;
    SS0[19][11] = 4'hE;
    SS0[20][11] = 4'hE;
    SS0[21][11] = 4'h0;
    SS0[22][11] = 4'h0;
    SS0[23][11] = 4'h0;
    SS0[24][11] = 4'h0;
    SS0[25][11] = 4'h0;
    SS0[26][11] = 4'h0;
    SS0[27][11] = 4'hE;
    SS0[28][11] = 4'hE;
    SS0[29][11] = 4'hE;
    SS0[30][11] = 4'hD;
    SS0[31][11] = 4'hD;
    SS0[32][11] = 4'hD;
    SS0[33][11] = 4'hC;
    SS0[34][11] = 4'hC;
    SS0[35][11] = 4'hC;
    SS0[36][11] = 4'h0;
    SS0[37][11] = 4'h0;
    SS0[38][11] = 4'h0;
    SS0[39][11] = 4'h0;
    SS0[40][11] = 4'h0;
    SS0[41][11] = 4'h0;
    SS0[42][11] = 4'h0;
    SS0[43][11] = 4'h0;
    SS0[44][11] = 4'h0;
    SS0[45][11] = 4'h0;
    SS0[46][11] = 4'h0;
    SS0[47][11] = 4'h0;
    SS0[0][12] = 4'h0;
    SS0[1][12] = 4'h0;
    SS0[2][12] = 4'h0;
    SS0[3][12] = 4'h0;
    SS0[4][12] = 4'h0;
    SS0[5][12] = 4'h0;
    SS0[6][12] = 4'h0;
    SS0[7][12] = 4'h0;
    SS0[8][12] = 4'h0;
    SS0[9][12] = 4'h0;
    SS0[10][12] = 4'h0;
    SS0[11][12] = 4'h0;
    SS0[12][12] = 4'hC;
    SS0[13][12] = 4'hC;
    SS0[14][12] = 4'hC;
    SS0[15][12] = 4'hC;
    SS0[16][12] = 4'hC;
    SS0[17][12] = 4'hC;
    SS0[18][12] = 4'hD;
    SS0[19][12] = 4'hD;
    SS0[20][12] = 4'hD;
    SS0[21][12] = 4'hE;
    SS0[22][12] = 4'hE;
    SS0[23][12] = 4'hE;
    SS0[24][12] = 4'hE;
    SS0[25][12] = 4'hE;
    SS0[26][12] = 4'hE;
    SS0[27][12] = 4'hD;
    SS0[28][12] = 4'hD;
    SS0[29][12] = 4'hD;
    SS0[30][12] = 4'hC;
    SS0[31][12] = 4'hC;
    SS0[32][12] = 4'hC;
    SS0[33][12] = 4'hC;
    SS0[34][12] = 4'hC;
    SS0[35][12] = 4'hC;
    SS0[36][12] = 4'h0;
    SS0[37][12] = 4'h0;
    SS0[38][12] = 4'h0;
    SS0[39][12] = 4'h0;
    SS0[40][12] = 4'h0;
    SS0[41][12] = 4'h0;
    SS0[42][12] = 4'h0;
    SS0[43][12] = 4'h0;
    SS0[44][12] = 4'h0;
    SS0[45][12] = 4'h0;
    SS0[46][12] = 4'h0;
    SS0[47][12] = 4'h0;
    SS0[0][13] = 4'h0;
    SS0[1][13] = 4'h0;
    SS0[2][13] = 4'h0;
    SS0[3][13] = 4'h0;
    SS0[4][13] = 4'h0;
    SS0[5][13] = 4'h0;
    SS0[6][13] = 4'h0;
    SS0[7][13] = 4'h0;
    SS0[8][13] = 4'h0;
    SS0[9][13] = 4'h0;
    SS0[10][13] = 4'h0;
    SS0[11][13] = 4'h0;
    SS0[12][13] = 4'hC;
    SS0[13][13] = 4'hC;
    SS0[14][13] = 4'hC;
    SS0[15][13] = 4'hC;
    SS0[16][13] = 4'hC;
    SS0[17][13] = 4'hC;
    SS0[18][13] = 4'hD;
    SS0[19][13] = 4'hD;
    SS0[20][13] = 4'hD;
    SS0[21][13] = 4'hE;
    SS0[22][13] = 4'hE;
    SS0[23][13] = 4'hE;
    SS0[24][13] = 4'hE;
    SS0[25][13] = 4'hE;
    SS0[26][13] = 4'hE;
    SS0[27][13] = 4'hD;
    SS0[28][13] = 4'hD;
    SS0[29][13] = 4'hD;
    SS0[30][13] = 4'hC;
    SS0[31][13] = 4'hC;
    SS0[32][13] = 4'hC;
    SS0[33][13] = 4'hC;
    SS0[34][13] = 4'hC;
    SS0[35][13] = 4'hC;
    SS0[36][13] = 4'h0;
    SS0[37][13] = 4'h0;
    SS0[38][13] = 4'h0;
    SS0[39][13] = 4'h0;
    SS0[40][13] = 4'h0;
    SS0[41][13] = 4'h0;
    SS0[42][13] = 4'h0;
    SS0[43][13] = 4'h0;
    SS0[44][13] = 4'h0;
    SS0[45][13] = 4'h0;
    SS0[46][13] = 4'h0;
    SS0[47][13] = 4'h0;
    SS0[0][14] = 4'h0;
    SS0[1][14] = 4'h0;
    SS0[2][14] = 4'h0;
    SS0[3][14] = 4'h0;
    SS0[4][14] = 4'h0;
    SS0[5][14] = 4'h0;
    SS0[6][14] = 4'h0;
    SS0[7][14] = 4'h0;
    SS0[8][14] = 4'h0;
    SS0[9][14] = 4'h0;
    SS0[10][14] = 4'h0;
    SS0[11][14] = 4'h0;
    SS0[12][14] = 4'hC;
    SS0[13][14] = 4'hC;
    SS0[14][14] = 4'hC;
    SS0[15][14] = 4'hC;
    SS0[16][14] = 4'hC;
    SS0[17][14] = 4'hC;
    SS0[18][14] = 4'hD;
    SS0[19][14] = 4'hD;
    SS0[20][14] = 4'hD;
    SS0[21][14] = 4'hE;
    SS0[22][14] = 4'hE;
    SS0[23][14] = 4'hE;
    SS0[24][14] = 4'hE;
    SS0[25][14] = 4'hE;
    SS0[26][14] = 4'hE;
    SS0[27][14] = 4'hD;
    SS0[28][14] = 4'hD;
    SS0[29][14] = 4'hD;
    SS0[30][14] = 4'hC;
    SS0[31][14] = 4'hC;
    SS0[32][14] = 4'hC;
    SS0[33][14] = 4'hC;
    SS0[34][14] = 4'hC;
    SS0[35][14] = 4'hC;
    SS0[36][14] = 4'h0;
    SS0[37][14] = 4'h0;
    SS0[38][14] = 4'h0;
    SS0[39][14] = 4'h0;
    SS0[40][14] = 4'h0;
    SS0[41][14] = 4'h0;
    SS0[42][14] = 4'h0;
    SS0[43][14] = 4'h0;
    SS0[44][14] = 4'h0;
    SS0[45][14] = 4'h0;
    SS0[46][14] = 4'h0;
    SS0[47][14] = 4'h0;
    SS0[0][15] = 4'hD;
    SS0[1][15] = 4'hD;
    SS0[2][15] = 4'hD;
    SS0[3][15] = 4'hD;
    SS0[4][15] = 4'hD;
    SS0[5][15] = 4'hD;
    SS0[6][15] = 4'hE;
    SS0[7][15] = 4'hE;
    SS0[8][15] = 4'hE;
    SS0[9][15] = 4'hE;
    SS0[10][15] = 4'hE;
    SS0[11][15] = 4'hE;
    SS0[12][15] = 4'hC;
    SS0[13][15] = 4'hC;
    SS0[14][15] = 4'hC;
    SS0[15][15] = 4'hC;
    SS0[16][15] = 4'hC;
    SS0[17][15] = 4'hC;
    SS0[18][15] = 4'hC;
    SS0[19][15] = 4'hC;
    SS0[20][15] = 4'hC;
    SS0[21][15] = 4'hE;
    SS0[22][15] = 4'hE;
    SS0[23][15] = 4'hE;
    SS0[24][15] = 4'hE;
    SS0[25][15] = 4'hE;
    SS0[26][15] = 4'hE;
    SS0[27][15] = 4'hC;
    SS0[28][15] = 4'hC;
    SS0[29][15] = 4'hC;
    SS0[30][15] = 4'hC;
    SS0[31][15] = 4'hC;
    SS0[32][15] = 4'hC;
    SS0[33][15] = 4'hC;
    SS0[34][15] = 4'hC;
    SS0[35][15] = 4'hC;
    SS0[36][15] = 4'hE;
    SS0[37][15] = 4'hE;
    SS0[38][15] = 4'hE;
    SS0[39][15] = 4'hE;
    SS0[40][15] = 4'hE;
    SS0[41][15] = 4'hE;
    SS0[42][15] = 4'hD;
    SS0[43][15] = 4'hD;
    SS0[44][15] = 4'hD;
    SS0[45][15] = 4'hD;
    SS0[46][15] = 4'hD;
    SS0[47][15] = 4'hD;
    SS0[0][16] = 4'hD;
    SS0[1][16] = 4'hD;
    SS0[2][16] = 4'hD;
    SS0[3][16] = 4'hD;
    SS0[4][16] = 4'hD;
    SS0[5][16] = 4'hD;
    SS0[6][16] = 4'hE;
    SS0[7][16] = 4'hE;
    SS0[8][16] = 4'hE;
    SS0[9][16] = 4'hE;
    SS0[10][16] = 4'hE;
    SS0[11][16] = 4'hE;
    SS0[12][16] = 4'hC;
    SS0[13][16] = 4'hC;
    SS0[14][16] = 4'hC;
    SS0[15][16] = 4'hC;
    SS0[16][16] = 4'hC;
    SS0[17][16] = 4'hC;
    SS0[18][16] = 4'hC;
    SS0[19][16] = 4'hC;
    SS0[20][16] = 4'hC;
    SS0[21][16] = 4'hE;
    SS0[22][16] = 4'hE;
    SS0[23][16] = 4'hE;
    SS0[24][16] = 4'hE;
    SS0[25][16] = 4'hE;
    SS0[26][16] = 4'hE;
    SS0[27][16] = 4'hC;
    SS0[28][16] = 4'hC;
    SS0[29][16] = 4'hC;
    SS0[30][16] = 4'hC;
    SS0[31][16] = 4'hC;
    SS0[32][16] = 4'hC;
    SS0[33][16] = 4'hC;
    SS0[34][16] = 4'hC;
    SS0[35][16] = 4'hC;
    SS0[36][16] = 4'hE;
    SS0[37][16] = 4'hE;
    SS0[38][16] = 4'hE;
    SS0[39][16] = 4'hE;
    SS0[40][16] = 4'hE;
    SS0[41][16] = 4'hE;
    SS0[42][16] = 4'hD;
    SS0[43][16] = 4'hD;
    SS0[44][16] = 4'hD;
    SS0[45][16] = 4'hD;
    SS0[46][16] = 4'hD;
    SS0[47][16] = 4'hD;
    SS0[0][17] = 4'hD;
    SS0[1][17] = 4'hD;
    SS0[2][17] = 4'hD;
    SS0[3][17] = 4'hD;
    SS0[4][17] = 4'hD;
    SS0[5][17] = 4'hD;
    SS0[6][17] = 4'hE;
    SS0[7][17] = 4'hE;
    SS0[8][17] = 4'hE;
    SS0[9][17] = 4'hE;
    SS0[10][17] = 4'hE;
    SS0[11][17] = 4'hE;
    SS0[12][17] = 4'hC;
    SS0[13][17] = 4'hC;
    SS0[14][17] = 4'hC;
    SS0[15][17] = 4'hC;
    SS0[16][17] = 4'hC;
    SS0[17][17] = 4'hC;
    SS0[18][17] = 4'hC;
    SS0[19][17] = 4'hC;
    SS0[20][17] = 4'hC;
    SS0[21][17] = 4'hE;
    SS0[22][17] = 4'hE;
    SS0[23][17] = 4'hE;
    SS0[24][17] = 4'hE;
    SS0[25][17] = 4'hE;
    SS0[26][17] = 4'hE;
    SS0[27][17] = 4'hC;
    SS0[28][17] = 4'hC;
    SS0[29][17] = 4'hC;
    SS0[30][17] = 4'hC;
    SS0[31][17] = 4'hC;
    SS0[32][17] = 4'hC;
    SS0[33][17] = 4'hC;
    SS0[34][17] = 4'hC;
    SS0[35][17] = 4'hC;
    SS0[36][17] = 4'hE;
    SS0[37][17] = 4'hE;
    SS0[38][17] = 4'hE;
    SS0[39][17] = 4'hE;
    SS0[40][17] = 4'hE;
    SS0[41][17] = 4'hE;
    SS0[42][17] = 4'hD;
    SS0[43][17] = 4'hD;
    SS0[44][17] = 4'hD;
    SS0[45][17] = 4'hD;
    SS0[46][17] = 4'hD;
    SS0[47][17] = 4'hD;
    SS0[0][18] = 4'h0;
    SS0[1][18] = 4'h0;
    SS0[2][18] = 4'h0;
    SS0[3][18] = 4'hD;
    SS0[4][18] = 4'hD;
    SS0[5][18] = 4'hD;
    SS0[6][18] = 4'hD;
    SS0[7][18] = 4'hD;
    SS0[8][18] = 4'hD;
    SS0[9][18] = 4'hE;
    SS0[10][18] = 4'hE;
    SS0[11][18] = 4'hE;
    SS0[12][18] = 4'hE;
    SS0[13][18] = 4'hE;
    SS0[14][18] = 4'hE;
    SS0[15][18] = 4'hC;
    SS0[16][18] = 4'hC;
    SS0[17][18] = 4'hC;
    SS0[18][18] = 4'hC;
    SS0[19][18] = 4'hC;
    SS0[20][18] = 4'hC;
    SS0[21][18] = 4'hD;
    SS0[22][18] = 4'hD;
    SS0[23][18] = 4'hD;
    SS0[24][18] = 4'hD;
    SS0[25][18] = 4'hD;
    SS0[26][18] = 4'hD;
    SS0[27][18] = 4'hC;
    SS0[28][18] = 4'hC;
    SS0[29][18] = 4'hC;
    SS0[30][18] = 4'hC;
    SS0[31][18] = 4'hC;
    SS0[32][18] = 4'hC;
    SS0[33][18] = 4'hE;
    SS0[34][18] = 4'hE;
    SS0[35][18] = 4'hE;
    SS0[36][18] = 4'hE;
    SS0[37][18] = 4'hE;
    SS0[38][18] = 4'hE;
    SS0[39][18] = 4'hD;
    SS0[40][18] = 4'hD;
    SS0[41][18] = 4'hD;
    SS0[42][18] = 4'hD;
    SS0[43][18] = 4'hD;
    SS0[44][18] = 4'hD;
    SS0[45][18] = 4'h0;
    SS0[46][18] = 4'h0;
    SS0[47][18] = 4'h0;
    SS0[0][19] = 4'h0;
    SS0[1][19] = 4'h0;
    SS0[2][19] = 4'h0;
    SS0[3][19] = 4'hD;
    SS0[4][19] = 4'hD;
    SS0[5][19] = 4'hD;
    SS0[6][19] = 4'hD;
    SS0[7][19] = 4'hD;
    SS0[8][19] = 4'hD;
    SS0[9][19] = 4'hE;
    SS0[10][19] = 4'hE;
    SS0[11][19] = 4'hE;
    SS0[12][19] = 4'hE;
    SS0[13][19] = 4'hE;
    SS0[14][19] = 4'hE;
    SS0[15][19] = 4'hC;
    SS0[16][19] = 4'hC;
    SS0[17][19] = 4'hC;
    SS0[18][19] = 4'hC;
    SS0[19][19] = 4'hC;
    SS0[20][19] = 4'hC;
    SS0[21][19] = 4'hD;
    SS0[22][19] = 4'hD;
    SS0[23][19] = 4'hD;
    SS0[24][19] = 4'hD;
    SS0[25][19] = 4'hD;
    SS0[26][19] = 4'hD;
    SS0[27][19] = 4'hC;
    SS0[28][19] = 4'hC;
    SS0[29][19] = 4'hC;
    SS0[30][19] = 4'hC;
    SS0[31][19] = 4'hC;
    SS0[32][19] = 4'hC;
    SS0[33][19] = 4'hE;
    SS0[34][19] = 4'hE;
    SS0[35][19] = 4'hE;
    SS0[36][19] = 4'hE;
    SS0[37][19] = 4'hE;
    SS0[38][19] = 4'hE;
    SS0[39][19] = 4'hD;
    SS0[40][19] = 4'hD;
    SS0[41][19] = 4'hD;
    SS0[42][19] = 4'hD;
    SS0[43][19] = 4'hD;
    SS0[44][19] = 4'hD;
    SS0[45][19] = 4'h0;
    SS0[46][19] = 4'h0;
    SS0[47][19] = 4'h0;
    SS0[0][20] = 4'h0;
    SS0[1][20] = 4'h0;
    SS0[2][20] = 4'h0;
    SS0[3][20] = 4'hD;
    SS0[4][20] = 4'hD;
    SS0[5][20] = 4'hD;
    SS0[6][20] = 4'hD;
    SS0[7][20] = 4'hD;
    SS0[8][20] = 4'hD;
    SS0[9][20] = 4'hE;
    SS0[10][20] = 4'hE;
    SS0[11][20] = 4'hE;
    SS0[12][20] = 4'hE;
    SS0[13][20] = 4'hE;
    SS0[14][20] = 4'hE;
    SS0[15][20] = 4'hC;
    SS0[16][20] = 4'hC;
    SS0[17][20] = 4'hC;
    SS0[18][20] = 4'hC;
    SS0[19][20] = 4'hC;
    SS0[20][20] = 4'hC;
    SS0[21][20] = 4'hD;
    SS0[22][20] = 4'hD;
    SS0[23][20] = 4'hD;
    SS0[24][20] = 4'hD;
    SS0[25][20] = 4'hD;
    SS0[26][20] = 4'hD;
    SS0[27][20] = 4'hC;
    SS0[28][20] = 4'hC;
    SS0[29][20] = 4'hC;
    SS0[30][20] = 4'hC;
    SS0[31][20] = 4'hC;
    SS0[32][20] = 4'hC;
    SS0[33][20] = 4'hE;
    SS0[34][20] = 4'hE;
    SS0[35][20] = 4'hE;
    SS0[36][20] = 4'hE;
    SS0[37][20] = 4'hE;
    SS0[38][20] = 4'hE;
    SS0[39][20] = 4'hD;
    SS0[40][20] = 4'hD;
    SS0[41][20] = 4'hD;
    SS0[42][20] = 4'hD;
    SS0[43][20] = 4'hD;
    SS0[44][20] = 4'hD;
    SS0[45][20] = 4'h0;
    SS0[46][20] = 4'h0;
    SS0[47][20] = 4'h0;
    SS0[0][21] = 4'h0;
    SS0[1][21] = 4'h0;
    SS0[2][21] = 4'h0;
    SS0[3][21] = 4'h0;
    SS0[4][21] = 4'h0;
    SS0[5][21] = 4'h0;
    SS0[6][21] = 4'h3;
    SS0[7][21] = 4'h3;
    SS0[8][21] = 4'h3;
    SS0[9][21] = 4'hD;
    SS0[10][21] = 4'hD;
    SS0[11][21] = 4'hD;
    SS0[12][21] = 4'hD;
    SS0[13][21] = 4'hD;
    SS0[14][21] = 4'hD;
    SS0[15][21] = 4'hE;
    SS0[16][21] = 4'hE;
    SS0[17][21] = 4'hE;
    SS0[18][21] = 4'hC;
    SS0[19][21] = 4'hC;
    SS0[20][21] = 4'hC;
    SS0[21][21] = 4'hC;
    SS0[22][21] = 4'hC;
    SS0[23][21] = 4'hC;
    SS0[24][21] = 4'hC;
    SS0[25][21] = 4'hC;
    SS0[26][21] = 4'hC;
    SS0[27][21] = 4'hC;
    SS0[28][21] = 4'hC;
    SS0[29][21] = 4'hC;
    SS0[30][21] = 4'hE;
    SS0[31][21] = 4'hE;
    SS0[32][21] = 4'hE;
    SS0[33][21] = 4'hD;
    SS0[34][21] = 4'hD;
    SS0[35][21] = 4'hD;
    SS0[36][21] = 4'hD;
    SS0[37][21] = 4'hD;
    SS0[38][21] = 4'hD;
    SS0[39][21] = 4'h3;
    SS0[40][21] = 4'h3;
    SS0[41][21] = 4'h3;
    SS0[42][21] = 4'h0;
    SS0[43][21] = 4'h0;
    SS0[44][21] = 4'h0;
    SS0[45][21] = 4'h0;
    SS0[46][21] = 4'h0;
    SS0[47][21] = 4'h0;
    SS0[0][22] = 4'h0;
    SS0[1][22] = 4'h0;
    SS0[2][22] = 4'h0;
    SS0[3][22] = 4'h0;
    SS0[4][22] = 4'h0;
    SS0[5][22] = 4'h0;
    SS0[6][22] = 4'h3;
    SS0[7][22] = 4'h3;
    SS0[8][22] = 4'h3;
    SS0[9][22] = 4'hD;
    SS0[10][22] = 4'hD;
    SS0[11][22] = 4'hD;
    SS0[12][22] = 4'hD;
    SS0[13][22] = 4'hD;
    SS0[14][22] = 4'hD;
    SS0[15][22] = 4'hE;
    SS0[16][22] = 4'hE;
    SS0[17][22] = 4'hE;
    SS0[18][22] = 4'hC;
    SS0[19][22] = 4'hC;
    SS0[20][22] = 4'hC;
    SS0[21][22] = 4'hC;
    SS0[22][22] = 4'hC;
    SS0[23][22] = 4'hC;
    SS0[24][22] = 4'hC;
    SS0[25][22] = 4'hC;
    SS0[26][22] = 4'hC;
    SS0[27][22] = 4'hC;
    SS0[28][22] = 4'hC;
    SS0[29][22] = 4'hC;
    SS0[30][22] = 4'hE;
    SS0[31][22] = 4'hE;
    SS0[32][22] = 4'hE;
    SS0[33][22] = 4'hD;
    SS0[34][22] = 4'hD;
    SS0[35][22] = 4'hD;
    SS0[36][22] = 4'hD;
    SS0[37][22] = 4'hD;
    SS0[38][22] = 4'hD;
    SS0[39][22] = 4'h3;
    SS0[40][22] = 4'h3;
    SS0[41][22] = 4'h3;
    SS0[42][22] = 4'h0;
    SS0[43][22] = 4'h0;
    SS0[44][22] = 4'h0;
    SS0[45][22] = 4'h0;
    SS0[46][22] = 4'h0;
    SS0[47][22] = 4'h0;
    SS0[0][23] = 4'h0;
    SS0[1][23] = 4'h0;
    SS0[2][23] = 4'h0;
    SS0[3][23] = 4'h0;
    SS0[4][23] = 4'h0;
    SS0[5][23] = 4'h0;
    SS0[6][23] = 4'h3;
    SS0[7][23] = 4'h3;
    SS0[8][23] = 4'h3;
    SS0[9][23] = 4'hD;
    SS0[10][23] = 4'hD;
    SS0[11][23] = 4'hD;
    SS0[12][23] = 4'hD;
    SS0[13][23] = 4'hD;
    SS0[14][23] = 4'hD;
    SS0[15][23] = 4'hE;
    SS0[16][23] = 4'hE;
    SS0[17][23] = 4'hE;
    SS0[18][23] = 4'hC;
    SS0[19][23] = 4'hC;
    SS0[20][23] = 4'hC;
    SS0[21][23] = 4'hC;
    SS0[22][23] = 4'hC;
    SS0[23][23] = 4'hC;
    SS0[24][23] = 4'hC;
    SS0[25][23] = 4'hC;
    SS0[26][23] = 4'hC;
    SS0[27][23] = 4'hC;
    SS0[28][23] = 4'hC;
    SS0[29][23] = 4'hC;
    SS0[30][23] = 4'hE;
    SS0[31][23] = 4'hE;
    SS0[32][23] = 4'hE;
    SS0[33][23] = 4'hD;
    SS0[34][23] = 4'hD;
    SS0[35][23] = 4'hD;
    SS0[36][23] = 4'hD;
    SS0[37][23] = 4'hD;
    SS0[38][23] = 4'hD;
    SS0[39][23] = 4'h3;
    SS0[40][23] = 4'h3;
    SS0[41][23] = 4'h3;
    SS0[42][23] = 4'h0;
    SS0[43][23] = 4'h0;
    SS0[44][23] = 4'h0;
    SS0[45][23] = 4'h0;
    SS0[46][23] = 4'h0;
    SS0[47][23] = 4'h0;
    SS0[0][24] = 4'h0;
    SS0[1][24] = 4'h0;
    SS0[2][24] = 4'h0;
    SS0[3][24] = 4'h0;
    SS0[4][24] = 4'h0;
    SS0[5][24] = 4'h0;
    SS0[6][24] = 4'h0;
    SS0[7][24] = 4'h0;
    SS0[8][24] = 4'h0;
    SS0[9][24] = 4'h0;
    SS0[10][24] = 4'h0;
    SS0[11][24] = 4'h0;
    SS0[12][24] = 4'hD;
    SS0[13][24] = 4'hD;
    SS0[14][24] = 4'hD;
    SS0[15][24] = 4'hD;
    SS0[16][24] = 4'hD;
    SS0[17][24] = 4'hD;
    SS0[18][24] = 4'hC;
    SS0[19][24] = 4'hC;
    SS0[20][24] = 4'hC;
    SS0[21][24] = 4'hD;
    SS0[22][24] = 4'hD;
    SS0[23][24] = 4'hD;
    SS0[24][24] = 4'hD;
    SS0[25][24] = 4'hD;
    SS0[26][24] = 4'hD;
    SS0[27][24] = 4'hC;
    SS0[28][24] = 4'hC;
    SS0[29][24] = 4'hC;
    SS0[30][24] = 4'hD;
    SS0[31][24] = 4'hD;
    SS0[32][24] = 4'hD;
    SS0[33][24] = 4'hD;
    SS0[34][24] = 4'hD;
    SS0[35][24] = 4'hD;
    SS0[36][24] = 4'h0;
    SS0[37][24] = 4'h0;
    SS0[38][24] = 4'h0;
    SS0[39][24] = 4'h0;
    SS0[40][24] = 4'h0;
    SS0[41][24] = 4'h0;
    SS0[42][24] = 4'h0;
    SS0[43][24] = 4'h0;
    SS0[44][24] = 4'h0;
    SS0[45][24] = 4'h0;
    SS0[46][24] = 4'h0;
    SS0[47][24] = 4'h0;
    SS0[0][25] = 4'h0;
    SS0[1][25] = 4'h0;
    SS0[2][25] = 4'h0;
    SS0[3][25] = 4'h0;
    SS0[4][25] = 4'h0;
    SS0[5][25] = 4'h0;
    SS0[6][25] = 4'h0;
    SS0[7][25] = 4'h0;
    SS0[8][25] = 4'h0;
    SS0[9][25] = 4'h0;
    SS0[10][25] = 4'h0;
    SS0[11][25] = 4'h0;
    SS0[12][25] = 4'hD;
    SS0[13][25] = 4'hD;
    SS0[14][25] = 4'hD;
    SS0[15][25] = 4'hD;
    SS0[16][25] = 4'hD;
    SS0[17][25] = 4'hD;
    SS0[18][25] = 4'hC;
    SS0[19][25] = 4'hC;
    SS0[20][25] = 4'hC;
    SS0[21][25] = 4'hD;
    SS0[22][25] = 4'hD;
    SS0[23][25] = 4'hD;
    SS0[24][25] = 4'hD;
    SS0[25][25] = 4'hD;
    SS0[26][25] = 4'hD;
    SS0[27][25] = 4'hC;
    SS0[28][25] = 4'hC;
    SS0[29][25] = 4'hC;
    SS0[30][25] = 4'hD;
    SS0[31][25] = 4'hD;
    SS0[32][25] = 4'hD;
    SS0[33][25] = 4'hD;
    SS0[34][25] = 4'hD;
    SS0[35][25] = 4'hD;
    SS0[36][25] = 4'h0;
    SS0[37][25] = 4'h0;
    SS0[38][25] = 4'h0;
    SS0[39][25] = 4'h0;
    SS0[40][25] = 4'h0;
    SS0[41][25] = 4'h0;
    SS0[42][25] = 4'h0;
    SS0[43][25] = 4'h0;
    SS0[44][25] = 4'h0;
    SS0[45][25] = 4'h0;
    SS0[46][25] = 4'h0;
    SS0[47][25] = 4'h0;
    SS0[0][26] = 4'h0;
    SS0[1][26] = 4'h0;
    SS0[2][26] = 4'h0;
    SS0[3][26] = 4'h0;
    SS0[4][26] = 4'h0;
    SS0[5][26] = 4'h0;
    SS0[6][26] = 4'h0;
    SS0[7][26] = 4'h0;
    SS0[8][26] = 4'h0;
    SS0[9][26] = 4'h0;
    SS0[10][26] = 4'h0;
    SS0[11][26] = 4'h0;
    SS0[12][26] = 4'hD;
    SS0[13][26] = 4'hD;
    SS0[14][26] = 4'hD;
    SS0[15][26] = 4'hD;
    SS0[16][26] = 4'hD;
    SS0[17][26] = 4'hD;
    SS0[18][26] = 4'hC;
    SS0[19][26] = 4'hC;
    SS0[20][26] = 4'hC;
    SS0[21][26] = 4'hD;
    SS0[22][26] = 4'hD;
    SS0[23][26] = 4'hD;
    SS0[24][26] = 4'hD;
    SS0[25][26] = 4'hD;
    SS0[26][26] = 4'hD;
    SS0[27][26] = 4'hC;
    SS0[28][26] = 4'hC;
    SS0[29][26] = 4'hC;
    SS0[30][26] = 4'hD;
    SS0[31][26] = 4'hD;
    SS0[32][26] = 4'hD;
    SS0[33][26] = 4'hD;
    SS0[34][26] = 4'hD;
    SS0[35][26] = 4'hD;
    SS0[36][26] = 4'h0;
    SS0[37][26] = 4'h0;
    SS0[38][26] = 4'h0;
    SS0[39][26] = 4'h0;
    SS0[40][26] = 4'h0;
    SS0[41][26] = 4'h0;
    SS0[42][26] = 4'h0;
    SS0[43][26] = 4'h0;
    SS0[44][26] = 4'h0;
    SS0[45][26] = 4'h0;
    SS0[46][26] = 4'h0;
    SS0[47][26] = 4'h0;
    SS0[0][27] = 4'h0;
    SS0[1][27] = 4'h0;
    SS0[2][27] = 4'h0;
    SS0[3][27] = 4'h0;
    SS0[4][27] = 4'h0;
    SS0[5][27] = 4'h0;
    SS0[6][27] = 4'h0;
    SS0[7][27] = 4'h0;
    SS0[8][27] = 4'h0;
    SS0[9][27] = 4'h0;
    SS0[10][27] = 4'h0;
    SS0[11][27] = 4'h0;
    SS0[12][27] = 4'h3;
    SS0[13][27] = 4'h3;
    SS0[14][27] = 4'h3;
    SS0[15][27] = 4'hD;
    SS0[16][27] = 4'hD;
    SS0[17][27] = 4'hD;
    SS0[18][27] = 4'hD;
    SS0[19][27] = 4'hD;
    SS0[20][27] = 4'hD;
    SS0[21][27] = 4'hA;
    SS0[22][27] = 4'hA;
    SS0[23][27] = 4'hA;
    SS0[24][27] = 4'hA;
    SS0[25][27] = 4'hA;
    SS0[26][27] = 4'hA;
    SS0[27][27] = 4'hD;
    SS0[28][27] = 4'hD;
    SS0[29][27] = 4'hD;
    SS0[30][27] = 4'hD;
    SS0[31][27] = 4'hD;
    SS0[32][27] = 4'hD;
    SS0[33][27] = 4'h3;
    SS0[34][27] = 4'h3;
    SS0[35][27] = 4'h3;
    SS0[36][27] = 4'h0;
    SS0[37][27] = 4'h0;
    SS0[38][27] = 4'h0;
    SS0[39][27] = 4'h0;
    SS0[40][27] = 4'h0;
    SS0[41][27] = 4'h0;
    SS0[42][27] = 4'h0;
    SS0[43][27] = 4'h0;
    SS0[44][27] = 4'h0;
    SS0[45][27] = 4'h0;
    SS0[46][27] = 4'h0;
    SS0[47][27] = 4'h0;
    SS0[0][28] = 4'h0;
    SS0[1][28] = 4'h0;
    SS0[2][28] = 4'h0;
    SS0[3][28] = 4'h0;
    SS0[4][28] = 4'h0;
    SS0[5][28] = 4'h0;
    SS0[6][28] = 4'h0;
    SS0[7][28] = 4'h0;
    SS0[8][28] = 4'h0;
    SS0[9][28] = 4'h0;
    SS0[10][28] = 4'h0;
    SS0[11][28] = 4'h0;
    SS0[12][28] = 4'h3;
    SS0[13][28] = 4'h3;
    SS0[14][28] = 4'h3;
    SS0[15][28] = 4'hD;
    SS0[16][28] = 4'hD;
    SS0[17][28] = 4'hD;
    SS0[18][28] = 4'hD;
    SS0[19][28] = 4'hD;
    SS0[20][28] = 4'hD;
    SS0[21][28] = 4'hA;
    SS0[22][28] = 4'hA;
    SS0[23][28] = 4'hA;
    SS0[24][28] = 4'hA;
    SS0[25][28] = 4'hA;
    SS0[26][28] = 4'hA;
    SS0[27][28] = 4'hD;
    SS0[28][28] = 4'hD;
    SS0[29][28] = 4'hD;
    SS0[30][28] = 4'hD;
    SS0[31][28] = 4'hD;
    SS0[32][28] = 4'hD;
    SS0[33][28] = 4'h3;
    SS0[34][28] = 4'h3;
    SS0[35][28] = 4'h3;
    SS0[36][28] = 4'h0;
    SS0[37][28] = 4'h0;
    SS0[38][28] = 4'h0;
    SS0[39][28] = 4'h0;
    SS0[40][28] = 4'h0;
    SS0[41][28] = 4'h0;
    SS0[42][28] = 4'h0;
    SS0[43][28] = 4'h0;
    SS0[44][28] = 4'h0;
    SS0[45][28] = 4'h0;
    SS0[46][28] = 4'h0;
    SS0[47][28] = 4'h0;
    SS0[0][29] = 4'h0;
    SS0[1][29] = 4'h0;
    SS0[2][29] = 4'h0;
    SS0[3][29] = 4'h0;
    SS0[4][29] = 4'h0;
    SS0[5][29] = 4'h0;
    SS0[6][29] = 4'h0;
    SS0[7][29] = 4'h0;
    SS0[8][29] = 4'h0;
    SS0[9][29] = 4'h0;
    SS0[10][29] = 4'h0;
    SS0[11][29] = 4'h0;
    SS0[12][29] = 4'h3;
    SS0[13][29] = 4'h3;
    SS0[14][29] = 4'h3;
    SS0[15][29] = 4'hD;
    SS0[16][29] = 4'hD;
    SS0[17][29] = 4'hD;
    SS0[18][29] = 4'hD;
    SS0[19][29] = 4'hD;
    SS0[20][29] = 4'hD;
    SS0[21][29] = 4'hA;
    SS0[22][29] = 4'hA;
    SS0[23][29] = 4'hA;
    SS0[24][29] = 4'hA;
    SS0[25][29] = 4'hA;
    SS0[26][29] = 4'hA;
    SS0[27][29] = 4'hD;
    SS0[28][29] = 4'hD;
    SS0[29][29] = 4'hD;
    SS0[30][29] = 4'hD;
    SS0[31][29] = 4'hD;
    SS0[32][29] = 4'hD;
    SS0[33][29] = 4'h3;
    SS0[34][29] = 4'h3;
    SS0[35][29] = 4'h3;
    SS0[36][29] = 4'h0;
    SS0[37][29] = 4'h0;
    SS0[38][29] = 4'h0;
    SS0[39][29] = 4'h0;
    SS0[40][29] = 4'h0;
    SS0[41][29] = 4'h0;
    SS0[42][29] = 4'h0;
    SS0[43][29] = 4'h0;
    SS0[44][29] = 4'h0;
    SS0[45][29] = 4'h0;
    SS0[46][29] = 4'h0;
    SS0[47][29] = 4'h0;
    SS0[0][30] = 4'h0;
    SS0[1][30] = 4'h0;
    SS0[2][30] = 4'h0;
    SS0[3][30] = 4'h0;
    SS0[4][30] = 4'h0;
    SS0[5][30] = 4'h0;
    SS0[6][30] = 4'h0;
    SS0[7][30] = 4'h0;
    SS0[8][30] = 4'h0;
    SS0[9][30] = 4'h0;
    SS0[10][30] = 4'h0;
    SS0[11][30] = 4'h0;
    SS0[12][30] = 4'h0;
    SS0[13][30] = 4'h0;
    SS0[14][30] = 4'h0;
    SS0[15][30] = 4'h0;
    SS0[16][30] = 4'h0;
    SS0[17][30] = 4'h0;
    SS0[18][30] = 4'hC;
    SS0[19][30] = 4'hC;
    SS0[20][30] = 4'hC;
    SS0[21][30] = 4'hC;
    SS0[22][30] = 4'hC;
    SS0[23][30] = 4'hC;
    SS0[24][30] = 4'hC;
    SS0[25][30] = 4'hC;
    SS0[26][30] = 4'hC;
    SS0[27][30] = 4'hC;
    SS0[28][30] = 4'hC;
    SS0[29][30] = 4'hC;
    SS0[30][30] = 4'h0;
    SS0[31][30] = 4'h0;
    SS0[32][30] = 4'h0;
    SS0[33][30] = 4'h0;
    SS0[34][30] = 4'h0;
    SS0[35][30] = 4'h0;
    SS0[36][30] = 4'h0;
    SS0[37][30] = 4'h0;
    SS0[38][30] = 4'h0;
    SS0[39][30] = 4'h0;
    SS0[40][30] = 4'h0;
    SS0[41][30] = 4'h0;
    SS0[42][30] = 4'h0;
    SS0[43][30] = 4'h0;
    SS0[44][30] = 4'h0;
    SS0[45][30] = 4'h0;
    SS0[46][30] = 4'h0;
    SS0[47][30] = 4'h0;
    SS0[0][31] = 4'h0;
    SS0[1][31] = 4'h0;
    SS0[2][31] = 4'h0;
    SS0[3][31] = 4'h0;
    SS0[4][31] = 4'h0;
    SS0[5][31] = 4'h0;
    SS0[6][31] = 4'h0;
    SS0[7][31] = 4'h0;
    SS0[8][31] = 4'h0;
    SS0[9][31] = 4'h0;
    SS0[10][31] = 4'h0;
    SS0[11][31] = 4'h0;
    SS0[12][31] = 4'h0;
    SS0[13][31] = 4'h0;
    SS0[14][31] = 4'h0;
    SS0[15][31] = 4'h0;
    SS0[16][31] = 4'h0;
    SS0[17][31] = 4'h0;
    SS0[18][31] = 4'hC;
    SS0[19][31] = 4'hC;
    SS0[20][31] = 4'hC;
    SS0[21][31] = 4'hC;
    SS0[22][31] = 4'hC;
    SS0[23][31] = 4'hC;
    SS0[24][31] = 4'hC;
    SS0[25][31] = 4'hC;
    SS0[26][31] = 4'hC;
    SS0[27][31] = 4'hC;
    SS0[28][31] = 4'hC;
    SS0[29][31] = 4'hC;
    SS0[30][31] = 4'h0;
    SS0[31][31] = 4'h0;
    SS0[32][31] = 4'h0;
    SS0[33][31] = 4'h0;
    SS0[34][31] = 4'h0;
    SS0[35][31] = 4'h0;
    SS0[36][31] = 4'h0;
    SS0[37][31] = 4'h0;
    SS0[38][31] = 4'h0;
    SS0[39][31] = 4'h0;
    SS0[40][31] = 4'h0;
    SS0[41][31] = 4'h0;
    SS0[42][31] = 4'h0;
    SS0[43][31] = 4'h0;
    SS0[44][31] = 4'h0;
    SS0[45][31] = 4'h0;
    SS0[46][31] = 4'h0;
    SS0[47][31] = 4'h0;
    SS0[0][32] = 4'h0;
    SS0[1][32] = 4'h0;
    SS0[2][32] = 4'h0;
    SS0[3][32] = 4'h0;
    SS0[4][32] = 4'h0;
    SS0[5][32] = 4'h0;
    SS0[6][32] = 4'h0;
    SS0[7][32] = 4'h0;
    SS0[8][32] = 4'h0;
    SS0[9][32] = 4'h0;
    SS0[10][32] = 4'h0;
    SS0[11][32] = 4'h0;
    SS0[12][32] = 4'h0;
    SS0[13][32] = 4'h0;
    SS0[14][32] = 4'h0;
    SS0[15][32] = 4'h0;
    SS0[16][32] = 4'h0;
    SS0[17][32] = 4'h0;
    SS0[18][32] = 4'hC;
    SS0[19][32] = 4'hC;
    SS0[20][32] = 4'hC;
    SS0[21][32] = 4'hC;
    SS0[22][32] = 4'hC;
    SS0[23][32] = 4'hC;
    SS0[24][32] = 4'hC;
    SS0[25][32] = 4'hC;
    SS0[26][32] = 4'hC;
    SS0[27][32] = 4'hC;
    SS0[28][32] = 4'hC;
    SS0[29][32] = 4'hC;
    SS0[30][32] = 4'h0;
    SS0[31][32] = 4'h0;
    SS0[32][32] = 4'h0;
    SS0[33][32] = 4'h0;
    SS0[34][32] = 4'h0;
    SS0[35][32] = 4'h0;
    SS0[36][32] = 4'h0;
    SS0[37][32] = 4'h0;
    SS0[38][32] = 4'h0;
    SS0[39][32] = 4'h0;
    SS0[40][32] = 4'h0;
    SS0[41][32] = 4'h0;
    SS0[42][32] = 4'h0;
    SS0[43][32] = 4'h0;
    SS0[44][32] = 4'h0;
    SS0[45][32] = 4'h0;
    SS0[46][32] = 4'h0;
    SS0[47][32] = 4'h0;
    SS0[0][33] = 4'h0;
    SS0[1][33] = 4'h0;
    SS0[2][33] = 4'h0;
    SS0[3][33] = 4'h0;
    SS0[4][33] = 4'h0;
    SS0[5][33] = 4'h0;
    SS0[6][33] = 4'h0;
    SS0[7][33] = 4'h0;
    SS0[8][33] = 4'h0;
    SS0[9][33] = 4'h0;
    SS0[10][33] = 4'h0;
    SS0[11][33] = 4'h0;
    SS0[12][33] = 4'h0;
    SS0[13][33] = 4'h0;
    SS0[14][33] = 4'h0;
    SS0[15][33] = 4'h0;
    SS0[16][33] = 4'h0;
    SS0[17][33] = 4'h0;
    SS0[18][33] = 4'hD;
    SS0[19][33] = 4'hD;
    SS0[20][33] = 4'hD;
    SS0[21][33] = 4'hC;
    SS0[22][33] = 4'hC;
    SS0[23][33] = 4'hC;
    SS0[24][33] = 4'hC;
    SS0[25][33] = 4'hC;
    SS0[26][33] = 4'hC;
    SS0[27][33] = 4'hD;
    SS0[28][33] = 4'hD;
    SS0[29][33] = 4'hD;
    SS0[30][33] = 4'h0;
    SS0[31][33] = 4'h0;
    SS0[32][33] = 4'h0;
    SS0[33][33] = 4'h0;
    SS0[34][33] = 4'h0;
    SS0[35][33] = 4'h0;
    SS0[36][33] = 4'h0;
    SS0[37][33] = 4'h0;
    SS0[38][33] = 4'h0;
    SS0[39][33] = 4'h0;
    SS0[40][33] = 4'h0;
    SS0[41][33] = 4'h0;
    SS0[42][33] = 4'h0;
    SS0[43][33] = 4'h0;
    SS0[44][33] = 4'h0;
    SS0[45][33] = 4'h0;
    SS0[46][33] = 4'h0;
    SS0[47][33] = 4'h0;
    SS0[0][34] = 4'h0;
    SS0[1][34] = 4'h0;
    SS0[2][34] = 4'h0;
    SS0[3][34] = 4'h0;
    SS0[4][34] = 4'h0;
    SS0[5][34] = 4'h0;
    SS0[6][34] = 4'h0;
    SS0[7][34] = 4'h0;
    SS0[8][34] = 4'h0;
    SS0[9][34] = 4'h0;
    SS0[10][34] = 4'h0;
    SS0[11][34] = 4'h0;
    SS0[12][34] = 4'h0;
    SS0[13][34] = 4'h0;
    SS0[14][34] = 4'h0;
    SS0[15][34] = 4'h0;
    SS0[16][34] = 4'h0;
    SS0[17][34] = 4'h0;
    SS0[18][34] = 4'hD;
    SS0[19][34] = 4'hD;
    SS0[20][34] = 4'hD;
    SS0[21][34] = 4'hC;
    SS0[22][34] = 4'hC;
    SS0[23][34] = 4'hC;
    SS0[24][34] = 4'hC;
    SS0[25][34] = 4'hC;
    SS0[26][34] = 4'hC;
    SS0[27][34] = 4'hD;
    SS0[28][34] = 4'hD;
    SS0[29][34] = 4'hD;
    SS0[30][34] = 4'h0;
    SS0[31][34] = 4'h0;
    SS0[32][34] = 4'h0;
    SS0[33][34] = 4'h0;
    SS0[34][34] = 4'h0;
    SS0[35][34] = 4'h0;
    SS0[36][34] = 4'h0;
    SS0[37][34] = 4'h0;
    SS0[38][34] = 4'h0;
    SS0[39][34] = 4'h0;
    SS0[40][34] = 4'h0;
    SS0[41][34] = 4'h0;
    SS0[42][34] = 4'h0;
    SS0[43][34] = 4'h0;
    SS0[44][34] = 4'h0;
    SS0[45][34] = 4'h0;
    SS0[46][34] = 4'h0;
    SS0[47][34] = 4'h0;
    SS0[0][35] = 4'h0;
    SS0[1][35] = 4'h0;
    SS0[2][35] = 4'h0;
    SS0[3][35] = 4'h0;
    SS0[4][35] = 4'h0;
    SS0[5][35] = 4'h0;
    SS0[6][35] = 4'h0;
    SS0[7][35] = 4'h0;
    SS0[8][35] = 4'h0;
    SS0[9][35] = 4'h0;
    SS0[10][35] = 4'h0;
    SS0[11][35] = 4'h0;
    SS0[12][35] = 4'h0;
    SS0[13][35] = 4'h0;
    SS0[14][35] = 4'h0;
    SS0[15][35] = 4'h0;
    SS0[16][35] = 4'h0;
    SS0[17][35] = 4'h0;
    SS0[18][35] = 4'hD;
    SS0[19][35] = 4'hD;
    SS0[20][35] = 4'hD;
    SS0[21][35] = 4'hC;
    SS0[22][35] = 4'hC;
    SS0[23][35] = 4'hC;
    SS0[24][35] = 4'hC;
    SS0[25][35] = 4'hC;
    SS0[26][35] = 4'hC;
    SS0[27][35] = 4'hD;
    SS0[28][35] = 4'hD;
    SS0[29][35] = 4'hD;
    SS0[30][35] = 4'h0;
    SS0[31][35] = 4'h0;
    SS0[32][35] = 4'h0;
    SS0[33][35] = 4'h0;
    SS0[34][35] = 4'h0;
    SS0[35][35] = 4'h0;
    SS0[36][35] = 4'h0;
    SS0[37][35] = 4'h0;
    SS0[38][35] = 4'h0;
    SS0[39][35] = 4'h0;
    SS0[40][35] = 4'h0;
    SS0[41][35] = 4'h0;
    SS0[42][35] = 4'h0;
    SS0[43][35] = 4'h0;
    SS0[44][35] = 4'h0;
    SS0[45][35] = 4'h0;
    SS0[46][35] = 4'h0;
    SS0[47][35] = 4'h0;
    SS0[0][36] = 4'h0;
    SS0[1][36] = 4'h0;
    SS0[2][36] = 4'h0;
    SS0[3][36] = 4'h0;
    SS0[4][36] = 4'h0;
    SS0[5][36] = 4'h0;
    SS0[6][36] = 4'h0;
    SS0[7][36] = 4'h0;
    SS0[8][36] = 4'h0;
    SS0[9][36] = 4'h0;
    SS0[10][36] = 4'h0;
    SS0[11][36] = 4'h0;
    SS0[12][36] = 4'h0;
    SS0[13][36] = 4'h0;
    SS0[14][36] = 4'h0;
    SS0[15][36] = 4'h0;
    SS0[16][36] = 4'h0;
    SS0[17][36] = 4'h0;
    SS0[18][36] = 4'hD;
    SS0[19][36] = 4'hD;
    SS0[20][36] = 4'hD;
    SS0[21][36] = 4'hC;
    SS0[22][36] = 4'hC;
    SS0[23][36] = 4'hC;
    SS0[24][36] = 4'hC;
    SS0[25][36] = 4'hC;
    SS0[26][36] = 4'hC;
    SS0[27][36] = 4'hD;
    SS0[28][36] = 4'hD;
    SS0[29][36] = 4'hD;
    SS0[30][36] = 4'h0;
    SS0[31][36] = 4'h0;
    SS0[32][36] = 4'h0;
    SS0[33][36] = 4'h0;
    SS0[34][36] = 4'h0;
    SS0[35][36] = 4'h0;
    SS0[36][36] = 4'h0;
    SS0[37][36] = 4'h0;
    SS0[38][36] = 4'h0;
    SS0[39][36] = 4'h0;
    SS0[40][36] = 4'h0;
    SS0[41][36] = 4'h0;
    SS0[42][36] = 4'h0;
    SS0[43][36] = 4'h0;
    SS0[44][36] = 4'h0;
    SS0[45][36] = 4'h0;
    SS0[46][36] = 4'h0;
    SS0[47][36] = 4'h0;
    SS0[0][37] = 4'h0;
    SS0[1][37] = 4'h0;
    SS0[2][37] = 4'h0;
    SS0[3][37] = 4'h0;
    SS0[4][37] = 4'h0;
    SS0[5][37] = 4'h0;
    SS0[6][37] = 4'h0;
    SS0[7][37] = 4'h0;
    SS0[8][37] = 4'h0;
    SS0[9][37] = 4'h0;
    SS0[10][37] = 4'h0;
    SS0[11][37] = 4'h0;
    SS0[12][37] = 4'h0;
    SS0[13][37] = 4'h0;
    SS0[14][37] = 4'h0;
    SS0[15][37] = 4'h0;
    SS0[16][37] = 4'h0;
    SS0[17][37] = 4'h0;
    SS0[18][37] = 4'hD;
    SS0[19][37] = 4'hD;
    SS0[20][37] = 4'hD;
    SS0[21][37] = 4'hC;
    SS0[22][37] = 4'hC;
    SS0[23][37] = 4'hC;
    SS0[24][37] = 4'hC;
    SS0[25][37] = 4'hC;
    SS0[26][37] = 4'hC;
    SS0[27][37] = 4'hD;
    SS0[28][37] = 4'hD;
    SS0[29][37] = 4'hD;
    SS0[30][37] = 4'h0;
    SS0[31][37] = 4'h0;
    SS0[32][37] = 4'h0;
    SS0[33][37] = 4'h0;
    SS0[34][37] = 4'h0;
    SS0[35][37] = 4'h0;
    SS0[36][37] = 4'h0;
    SS0[37][37] = 4'h0;
    SS0[38][37] = 4'h0;
    SS0[39][37] = 4'h0;
    SS0[40][37] = 4'h0;
    SS0[41][37] = 4'h0;
    SS0[42][37] = 4'h0;
    SS0[43][37] = 4'h0;
    SS0[44][37] = 4'h0;
    SS0[45][37] = 4'h0;
    SS0[46][37] = 4'h0;
    SS0[47][37] = 4'h0;
    SS0[0][38] = 4'h0;
    SS0[1][38] = 4'h0;
    SS0[2][38] = 4'h0;
    SS0[3][38] = 4'h0;
    SS0[4][38] = 4'h0;
    SS0[5][38] = 4'h0;
    SS0[6][38] = 4'h0;
    SS0[7][38] = 4'h0;
    SS0[8][38] = 4'h0;
    SS0[9][38] = 4'h0;
    SS0[10][38] = 4'h0;
    SS0[11][38] = 4'h0;
    SS0[12][38] = 4'h0;
    SS0[13][38] = 4'h0;
    SS0[14][38] = 4'h0;
    SS0[15][38] = 4'h0;
    SS0[16][38] = 4'h0;
    SS0[17][38] = 4'h0;
    SS0[18][38] = 4'hD;
    SS0[19][38] = 4'hD;
    SS0[20][38] = 4'hD;
    SS0[21][38] = 4'hC;
    SS0[22][38] = 4'hC;
    SS0[23][38] = 4'hC;
    SS0[24][38] = 4'hC;
    SS0[25][38] = 4'hC;
    SS0[26][38] = 4'hC;
    SS0[27][38] = 4'hD;
    SS0[28][38] = 4'hD;
    SS0[29][38] = 4'hD;
    SS0[30][38] = 4'h0;
    SS0[31][38] = 4'h0;
    SS0[32][38] = 4'h0;
    SS0[33][38] = 4'h0;
    SS0[34][38] = 4'h0;
    SS0[35][38] = 4'h0;
    SS0[36][38] = 4'h0;
    SS0[37][38] = 4'h0;
    SS0[38][38] = 4'h0;
    SS0[39][38] = 4'h0;
    SS0[40][38] = 4'h0;
    SS0[41][38] = 4'h0;
    SS0[42][38] = 4'h0;
    SS0[43][38] = 4'h0;
    SS0[44][38] = 4'h0;
    SS0[45][38] = 4'h0;
    SS0[46][38] = 4'h0;
    SS0[47][38] = 4'h0;
    SS0[0][39] = 4'h0;
    SS0[1][39] = 4'h0;
    SS0[2][39] = 4'h0;
    SS0[3][39] = 4'h0;
    SS0[4][39] = 4'h0;
    SS0[5][39] = 4'h0;
    SS0[6][39] = 4'h0;
    SS0[7][39] = 4'h0;
    SS0[8][39] = 4'h0;
    SS0[9][39] = 4'h0;
    SS0[10][39] = 4'h0;
    SS0[11][39] = 4'h0;
    SS0[12][39] = 4'h0;
    SS0[13][39] = 4'h0;
    SS0[14][39] = 4'h0;
    SS0[15][39] = 4'h0;
    SS0[16][39] = 4'h0;
    SS0[17][39] = 4'h0;
    SS0[18][39] = 4'hD;
    SS0[19][39] = 4'hD;
    SS0[20][39] = 4'hD;
    SS0[21][39] = 4'hC;
    SS0[22][39] = 4'hC;
    SS0[23][39] = 4'hC;
    SS0[24][39] = 4'hC;
    SS0[25][39] = 4'hC;
    SS0[26][39] = 4'hC;
    SS0[27][39] = 4'hD;
    SS0[28][39] = 4'hD;
    SS0[29][39] = 4'hD;
    SS0[30][39] = 4'h0;
    SS0[31][39] = 4'h0;
    SS0[32][39] = 4'h0;
    SS0[33][39] = 4'h0;
    SS0[34][39] = 4'h0;
    SS0[35][39] = 4'h0;
    SS0[36][39] = 4'h0;
    SS0[37][39] = 4'h0;
    SS0[38][39] = 4'h0;
    SS0[39][39] = 4'h0;
    SS0[40][39] = 4'h0;
    SS0[41][39] = 4'h0;
    SS0[42][39] = 4'h0;
    SS0[43][39] = 4'h0;
    SS0[44][39] = 4'h0;
    SS0[45][39] = 4'h0;
    SS0[46][39] = 4'h0;
    SS0[47][39] = 4'h0;
    SS0[0][40] = 4'h0;
    SS0[1][40] = 4'h0;
    SS0[2][40] = 4'h0;
    SS0[3][40] = 4'h0;
    SS0[4][40] = 4'h0;
    SS0[5][40] = 4'h0;
    SS0[6][40] = 4'h0;
    SS0[7][40] = 4'h0;
    SS0[8][40] = 4'h0;
    SS0[9][40] = 4'h0;
    SS0[10][40] = 4'h0;
    SS0[11][40] = 4'h0;
    SS0[12][40] = 4'h0;
    SS0[13][40] = 4'h0;
    SS0[14][40] = 4'h0;
    SS0[15][40] = 4'h0;
    SS0[16][40] = 4'h0;
    SS0[17][40] = 4'h0;
    SS0[18][40] = 4'hD;
    SS0[19][40] = 4'hD;
    SS0[20][40] = 4'hD;
    SS0[21][40] = 4'hC;
    SS0[22][40] = 4'hC;
    SS0[23][40] = 4'hC;
    SS0[24][40] = 4'hC;
    SS0[25][40] = 4'hC;
    SS0[26][40] = 4'hC;
    SS0[27][40] = 4'hD;
    SS0[28][40] = 4'hD;
    SS0[29][40] = 4'hD;
    SS0[30][40] = 4'h0;
    SS0[31][40] = 4'h0;
    SS0[32][40] = 4'h0;
    SS0[33][40] = 4'h0;
    SS0[34][40] = 4'h0;
    SS0[35][40] = 4'h0;
    SS0[36][40] = 4'h0;
    SS0[37][40] = 4'h0;
    SS0[38][40] = 4'h0;
    SS0[39][40] = 4'h0;
    SS0[40][40] = 4'h0;
    SS0[41][40] = 4'h0;
    SS0[42][40] = 4'h0;
    SS0[43][40] = 4'h0;
    SS0[44][40] = 4'h0;
    SS0[45][40] = 4'h0;
    SS0[46][40] = 4'h0;
    SS0[47][40] = 4'h0;
    SS0[0][41] = 4'h0;
    SS0[1][41] = 4'h0;
    SS0[2][41] = 4'h0;
    SS0[3][41] = 4'h0;
    SS0[4][41] = 4'h0;
    SS0[5][41] = 4'h0;
    SS0[6][41] = 4'h0;
    SS0[7][41] = 4'h0;
    SS0[8][41] = 4'h0;
    SS0[9][41] = 4'h0;
    SS0[10][41] = 4'h0;
    SS0[11][41] = 4'h0;
    SS0[12][41] = 4'h0;
    SS0[13][41] = 4'h0;
    SS0[14][41] = 4'h0;
    SS0[15][41] = 4'h0;
    SS0[16][41] = 4'h0;
    SS0[17][41] = 4'h0;
    SS0[18][41] = 4'hD;
    SS0[19][41] = 4'hD;
    SS0[20][41] = 4'hD;
    SS0[21][41] = 4'hC;
    SS0[22][41] = 4'hC;
    SS0[23][41] = 4'hC;
    SS0[24][41] = 4'hC;
    SS0[25][41] = 4'hC;
    SS0[26][41] = 4'hC;
    SS0[27][41] = 4'hD;
    SS0[28][41] = 4'hD;
    SS0[29][41] = 4'hD;
    SS0[30][41] = 4'h0;
    SS0[31][41] = 4'h0;
    SS0[32][41] = 4'h0;
    SS0[33][41] = 4'h0;
    SS0[34][41] = 4'h0;
    SS0[35][41] = 4'h0;
    SS0[36][41] = 4'h0;
    SS0[37][41] = 4'h0;
    SS0[38][41] = 4'h0;
    SS0[39][41] = 4'h0;
    SS0[40][41] = 4'h0;
    SS0[41][41] = 4'h0;
    SS0[42][41] = 4'h0;
    SS0[43][41] = 4'h0;
    SS0[44][41] = 4'h0;
    SS0[45][41] = 4'h0;
    SS0[46][41] = 4'h0;
    SS0[47][41] = 4'h0;
    SS0[0][42] = 4'h0;
    SS0[1][42] = 4'h0;
    SS0[2][42] = 4'h0;
    SS0[3][42] = 4'h0;
    SS0[4][42] = 4'h0;
    SS0[5][42] = 4'h0;
    SS0[6][42] = 4'h0;
    SS0[7][42] = 4'h0;
    SS0[8][42] = 4'h0;
    SS0[9][42] = 4'h0;
    SS0[10][42] = 4'h0;
    SS0[11][42] = 4'h0;
    SS0[12][42] = 4'h0;
    SS0[13][42] = 4'h0;
    SS0[14][42] = 4'h0;
    SS0[15][42] = 4'h0;
    SS0[16][42] = 4'h0;
    SS0[17][42] = 4'h0;
    SS0[18][42] = 4'h0;
    SS0[19][42] = 4'h0;
    SS0[20][42] = 4'h0;
    SS0[21][42] = 4'hC;
    SS0[22][42] = 4'hC;
    SS0[23][42] = 4'hC;
    SS0[24][42] = 4'hC;
    SS0[25][42] = 4'hC;
    SS0[26][42] = 4'hC;
    SS0[27][42] = 4'h0;
    SS0[28][42] = 4'h0;
    SS0[29][42] = 4'h0;
    SS0[30][42] = 4'h0;
    SS0[31][42] = 4'h0;
    SS0[32][42] = 4'h0;
    SS0[33][42] = 4'h0;
    SS0[34][42] = 4'h0;
    SS0[35][42] = 4'h0;
    SS0[36][42] = 4'h0;
    SS0[37][42] = 4'h0;
    SS0[38][42] = 4'h0;
    SS0[39][42] = 4'h0;
    SS0[40][42] = 4'h0;
    SS0[41][42] = 4'h0;
    SS0[42][42] = 4'h0;
    SS0[43][42] = 4'h0;
    SS0[44][42] = 4'h0;
    SS0[45][42] = 4'h0;
    SS0[46][42] = 4'h0;
    SS0[47][42] = 4'h0;
    SS0[0][43] = 4'h0;
    SS0[1][43] = 4'h0;
    SS0[2][43] = 4'h0;
    SS0[3][43] = 4'h0;
    SS0[4][43] = 4'h0;
    SS0[5][43] = 4'h0;
    SS0[6][43] = 4'h0;
    SS0[7][43] = 4'h0;
    SS0[8][43] = 4'h0;
    SS0[9][43] = 4'h0;
    SS0[10][43] = 4'h0;
    SS0[11][43] = 4'h0;
    SS0[12][43] = 4'h0;
    SS0[13][43] = 4'h0;
    SS0[14][43] = 4'h0;
    SS0[15][43] = 4'h0;
    SS0[16][43] = 4'h0;
    SS0[17][43] = 4'h0;
    SS0[18][43] = 4'h0;
    SS0[19][43] = 4'h0;
    SS0[20][43] = 4'h0;
    SS0[21][43] = 4'hC;
    SS0[22][43] = 4'hC;
    SS0[23][43] = 4'hC;
    SS0[24][43] = 4'hC;
    SS0[25][43] = 4'hC;
    SS0[26][43] = 4'hC;
    SS0[27][43] = 4'h0;
    SS0[28][43] = 4'h0;
    SS0[29][43] = 4'h0;
    SS0[30][43] = 4'h0;
    SS0[31][43] = 4'h0;
    SS0[32][43] = 4'h0;
    SS0[33][43] = 4'h0;
    SS0[34][43] = 4'h0;
    SS0[35][43] = 4'h0;
    SS0[36][43] = 4'h0;
    SS0[37][43] = 4'h0;
    SS0[38][43] = 4'h0;
    SS0[39][43] = 4'h0;
    SS0[40][43] = 4'h0;
    SS0[41][43] = 4'h0;
    SS0[42][43] = 4'h0;
    SS0[43][43] = 4'h0;
    SS0[44][43] = 4'h0;
    SS0[45][43] = 4'h0;
    SS0[46][43] = 4'h0;
    SS0[47][43] = 4'h0;
    SS0[0][44] = 4'h0;
    SS0[1][44] = 4'h0;
    SS0[2][44] = 4'h0;
    SS0[3][44] = 4'h0;
    SS0[4][44] = 4'h0;
    SS0[5][44] = 4'h0;
    SS0[6][44] = 4'h0;
    SS0[7][44] = 4'h0;
    SS0[8][44] = 4'h0;
    SS0[9][44] = 4'h0;
    SS0[10][44] = 4'h0;
    SS0[11][44] = 4'h0;
    SS0[12][44] = 4'h0;
    SS0[13][44] = 4'h0;
    SS0[14][44] = 4'h0;
    SS0[15][44] = 4'h0;
    SS0[16][44] = 4'h0;
    SS0[17][44] = 4'h0;
    SS0[18][44] = 4'h0;
    SS0[19][44] = 4'h0;
    SS0[20][44] = 4'h0;
    SS0[21][44] = 4'hC;
    SS0[22][44] = 4'hC;
    SS0[23][44] = 4'hC;
    SS0[24][44] = 4'hC;
    SS0[25][44] = 4'hC;
    SS0[26][44] = 4'hC;
    SS0[27][44] = 4'h0;
    SS0[28][44] = 4'h0;
    SS0[29][44] = 4'h0;
    SS0[30][44] = 4'h0;
    SS0[31][44] = 4'h0;
    SS0[32][44] = 4'h0;
    SS0[33][44] = 4'h0;
    SS0[34][44] = 4'h0;
    SS0[35][44] = 4'h0;
    SS0[36][44] = 4'h0;
    SS0[37][44] = 4'h0;
    SS0[38][44] = 4'h0;
    SS0[39][44] = 4'h0;
    SS0[40][44] = 4'h0;
    SS0[41][44] = 4'h0;
    SS0[42][44] = 4'h0;
    SS0[43][44] = 4'h0;
    SS0[44][44] = 4'h0;
    SS0[45][44] = 4'h0;
    SS0[46][44] = 4'h0;
    SS0[47][44] = 4'h0;
    SS0[0][45] = 4'h0;
    SS0[1][45] = 4'h0;
    SS0[2][45] = 4'h0;
    SS0[3][45] = 4'h0;
    SS0[4][45] = 4'h0;
    SS0[5][45] = 4'h0;
    SS0[6][45] = 4'h0;
    SS0[7][45] = 4'h0;
    SS0[8][45] = 4'h0;
    SS0[9][45] = 4'h0;
    SS0[10][45] = 4'h0;
    SS0[11][45] = 4'h0;
    SS0[12][45] = 4'h0;
    SS0[13][45] = 4'h0;
    SS0[14][45] = 4'h0;
    SS0[15][45] = 4'h0;
    SS0[16][45] = 4'h0;
    SS0[17][45] = 4'h0;
    SS0[18][45] = 4'h0;
    SS0[19][45] = 4'h0;
    SS0[20][45] = 4'h0;
    SS0[21][45] = 4'hC;
    SS0[22][45] = 4'hC;
    SS0[23][45] = 4'hC;
    SS0[24][45] = 4'hC;
    SS0[25][45] = 4'hC;
    SS0[26][45] = 4'hC;
    SS0[27][45] = 4'h0;
    SS0[28][45] = 4'h0;
    SS0[29][45] = 4'h0;
    SS0[30][45] = 4'h0;
    SS0[31][45] = 4'h0;
    SS0[32][45] = 4'h0;
    SS0[33][45] = 4'h0;
    SS0[34][45] = 4'h0;
    SS0[35][45] = 4'h0;
    SS0[36][45] = 4'h0;
    SS0[37][45] = 4'h0;
    SS0[38][45] = 4'h0;
    SS0[39][45] = 4'h0;
    SS0[40][45] = 4'h0;
    SS0[41][45] = 4'h0;
    SS0[42][45] = 4'h0;
    SS0[43][45] = 4'h0;
    SS0[44][45] = 4'h0;
    SS0[45][45] = 4'h0;
    SS0[46][45] = 4'h0;
    SS0[47][45] = 4'h0;
    SS0[0][46] = 4'h0;
    SS0[1][46] = 4'h0;
    SS0[2][46] = 4'h0;
    SS0[3][46] = 4'h0;
    SS0[4][46] = 4'h0;
    SS0[5][46] = 4'h0;
    SS0[6][46] = 4'h0;
    SS0[7][46] = 4'h0;
    SS0[8][46] = 4'h0;
    SS0[9][46] = 4'h0;
    SS0[10][46] = 4'h0;
    SS0[11][46] = 4'h0;
    SS0[12][46] = 4'h0;
    SS0[13][46] = 4'h0;
    SS0[14][46] = 4'h0;
    SS0[15][46] = 4'h0;
    SS0[16][46] = 4'h0;
    SS0[17][46] = 4'h0;
    SS0[18][46] = 4'h0;
    SS0[19][46] = 4'h0;
    SS0[20][46] = 4'h0;
    SS0[21][46] = 4'hC;
    SS0[22][46] = 4'hC;
    SS0[23][46] = 4'hC;
    SS0[24][46] = 4'hC;
    SS0[25][46] = 4'hC;
    SS0[26][46] = 4'hC;
    SS0[27][46] = 4'h0;
    SS0[28][46] = 4'h0;
    SS0[29][46] = 4'h0;
    SS0[30][46] = 4'h0;
    SS0[31][46] = 4'h0;
    SS0[32][46] = 4'h0;
    SS0[33][46] = 4'h0;
    SS0[34][46] = 4'h0;
    SS0[35][46] = 4'h0;
    SS0[36][46] = 4'h0;
    SS0[37][46] = 4'h0;
    SS0[38][46] = 4'h0;
    SS0[39][46] = 4'h0;
    SS0[40][46] = 4'h0;
    SS0[41][46] = 4'h0;
    SS0[42][46] = 4'h0;
    SS0[43][46] = 4'h0;
    SS0[44][46] = 4'h0;
    SS0[45][46] = 4'h0;
    SS0[46][46] = 4'h0;
    SS0[47][46] = 4'h0;
    SS0[0][47] = 4'h0;
    SS0[1][47] = 4'h0;
    SS0[2][47] = 4'h0;
    SS0[3][47] = 4'h0;
    SS0[4][47] = 4'h0;
    SS0[5][47] = 4'h0;
    SS0[6][47] = 4'h0;
    SS0[7][47] = 4'h0;
    SS0[8][47] = 4'h0;
    SS0[9][47] = 4'h0;
    SS0[10][47] = 4'h0;
    SS0[11][47] = 4'h0;
    SS0[12][47] = 4'h0;
    SS0[13][47] = 4'h0;
    SS0[14][47] = 4'h0;
    SS0[15][47] = 4'h0;
    SS0[16][47] = 4'h0;
    SS0[17][47] = 4'h0;
    SS0[18][47] = 4'h0;
    SS0[19][47] = 4'h0;
    SS0[20][47] = 4'h0;
    SS0[21][47] = 4'hC;
    SS0[22][47] = 4'hC;
    SS0[23][47] = 4'hC;
    SS0[24][47] = 4'hC;
    SS0[25][47] = 4'hC;
    SS0[26][47] = 4'hC;
    SS0[27][47] = 4'h0;
    SS0[28][47] = 4'h0;
    SS0[29][47] = 4'h0;
    SS0[30][47] = 4'h0;
    SS0[31][47] = 4'h0;
    SS0[32][47] = 4'h0;
    SS0[33][47] = 4'h0;
    SS0[34][47] = 4'h0;
    SS0[35][47] = 4'h0;
    SS0[36][47] = 4'h0;
    SS0[37][47] = 4'h0;
    SS0[38][47] = 4'h0;
    SS0[39][47] = 4'h0;
    SS0[40][47] = 4'h0;
    SS0[41][47] = 4'h0;
    SS0[42][47] = 4'h0;
    SS0[43][47] = 4'h0;
    SS0[44][47] = 4'h0;
    SS0[45][47] = 4'h0;
    SS0[46][47] = 4'h0;
    SS0[47][47] = 4'h0;
 
//SS 1
    SS1[0][0] = 4'h0;
    SS1[1][0] = 4'h0;
    SS1[2][0] = 4'h0;
    SS1[3][0] = 4'h0;
    SS1[4][0] = 4'h0;
    SS1[5][0] = 4'h0;
    SS1[6][0] = 4'h0;
    SS1[7][0] = 4'h0;
    SS1[8][0] = 4'h0;
    SS1[9][0] = 4'h0;
    SS1[10][0] = 4'h0;
    SS1[11][0] = 4'h0;
    SS1[12][0] = 4'h0;
    SS1[13][0] = 4'h0;
    SS1[14][0] = 4'h0;
    SS1[15][0] = 4'h0;
    SS1[16][0] = 4'h0;
    SS1[17][0] = 4'h0;
    SS1[18][0] = 4'hC;
    SS1[19][0] = 4'hC;
    SS1[20][0] = 4'hC;
    SS1[21][0] = 4'h0;
    SS1[22][0] = 4'h0;
    SS1[23][0] = 4'h0;
    SS1[24][0] = 4'h0;
    SS1[25][0] = 4'h0;
    SS1[26][0] = 4'h0;
    SS1[27][0] = 4'h0;
    SS1[28][0] = 4'h0;
    SS1[29][0] = 4'h0;
    SS1[30][0] = 4'h0;
    SS1[31][0] = 4'h0;
    SS1[32][0] = 4'h0;
    SS1[33][0] = 4'h0;
    SS1[34][0] = 4'h0;
    SS1[35][0] = 4'h0;
    SS1[36][0] = 4'h0;
    SS1[37][0] = 4'h0;
    SS1[38][0] = 4'h0;
    SS1[39][0] = 4'h0;
    SS1[40][0] = 4'h0;
    SS1[41][0] = 4'h0;
    SS1[42][0] = 4'h0;
    SS1[43][0] = 4'h0;
    SS1[44][0] = 4'h0;
    SS1[45][0] = 4'h0;
    SS1[46][0] = 4'h0;
    SS1[47][0] = 4'h0;
    SS1[0][1] = 4'h0;
    SS1[1][1] = 4'h0;
    SS1[2][1] = 4'h0;
    SS1[3][1] = 4'h0;
    SS1[4][1] = 4'h0;
    SS1[5][1] = 4'h0;
    SS1[6][1] = 4'h0;
    SS1[7][1] = 4'h0;
    SS1[8][1] = 4'h0;
    SS1[9][1] = 4'h0;
    SS1[10][1] = 4'h0;
    SS1[11][1] = 4'h0;
    SS1[12][1] = 4'h0;
    SS1[13][1] = 4'h0;
    SS1[14][1] = 4'h0;
    SS1[15][1] = 4'h0;
    SS1[16][1] = 4'h0;
    SS1[17][1] = 4'hC;
    SS1[18][1] = 4'hC;
    SS1[19][1] = 4'hC;
    SS1[20][1] = 4'hD;
    SS1[21][1] = 4'hD;
    SS1[22][1] = 4'hD;
    SS1[23][1] = 4'hD;
    SS1[24][1] = 4'h0;
    SS1[25][1] = 4'h0;
    SS1[26][1] = 4'h0;
    SS1[27][1] = 4'h0;
    SS1[28][1] = 4'h0;
    SS1[29][1] = 4'h0;
    SS1[30][1] = 4'h0;
    SS1[31][1] = 4'h0;
    SS1[32][1] = 4'h0;
    SS1[33][1] = 4'h0;
    SS1[34][1] = 4'h0;
    SS1[35][1] = 4'h0;
    SS1[36][1] = 4'h0;
    SS1[37][1] = 4'h0;
    SS1[38][1] = 4'h0;
    SS1[39][1] = 4'h0;
    SS1[40][1] = 4'h0;
    SS1[41][1] = 4'h0;
    SS1[42][1] = 4'h0;
    SS1[43][1] = 4'h0;
    SS1[44][1] = 4'h0;
    SS1[45][1] = 4'h0;
    SS1[46][1] = 4'h0;
    SS1[47][1] = 4'h0;
    SS1[0][2] = 4'h0;
    SS1[1][2] = 4'h0;
    SS1[2][2] = 4'h0;
    SS1[3][2] = 4'h0;
    SS1[4][2] = 4'h0;
    SS1[5][2] = 4'h0;
    SS1[6][2] = 4'h0;
    SS1[7][2] = 4'h0;
    SS1[8][2] = 4'h0;
    SS1[9][2] = 4'h0;
    SS1[10][2] = 4'h0;
    SS1[11][2] = 4'h0;
    SS1[12][2] = 4'h0;
    SS1[13][2] = 4'h0;
    SS1[14][2] = 4'h0;
    SS1[15][2] = 4'h0;
    SS1[16][2] = 4'h0;
    SS1[17][2] = 4'hC;
    SS1[18][2] = 4'hC;
    SS1[19][2] = 4'hC;
    SS1[20][2] = 4'hD;
    SS1[21][2] = 4'hD;
    SS1[22][2] = 4'hD;
    SS1[23][2] = 4'h0;
    SS1[24][2] = 4'h0;
    SS1[25][2] = 4'h0;
    SS1[26][2] = 4'h0;
    SS1[27][2] = 4'h0;
    SS1[28][2] = 4'h0;
    SS1[29][2] = 4'h0;
    SS1[30][2] = 4'h0;
    SS1[31][2] = 4'h0;
    SS1[32][2] = 4'h0;
    SS1[33][2] = 4'h0;
    SS1[34][2] = 4'h0;
    SS1[35][2] = 4'h0;
    SS1[36][2] = 4'h0;
    SS1[37][2] = 4'h0;
    SS1[38][2] = 4'h0;
    SS1[39][2] = 4'h0;
    SS1[40][2] = 4'h0;
    SS1[41][2] = 4'h0;
    SS1[42][2] = 4'h0;
    SS1[43][2] = 4'h0;
    SS1[44][2] = 4'h0;
    SS1[45][2] = 4'h0;
    SS1[46][2] = 4'h0;
    SS1[47][2] = 4'h0;
    SS1[0][3] = 4'h0;
    SS1[1][3] = 4'h0;
    SS1[2][3] = 4'h0;
    SS1[3][3] = 4'h0;
    SS1[4][3] = 4'h0;
    SS1[5][3] = 4'h0;
    SS1[6][3] = 4'h0;
    SS1[7][3] = 4'h0;
    SS1[8][3] = 4'h0;
    SS1[9][3] = 4'h0;
    SS1[10][3] = 4'h0;
    SS1[11][3] = 4'h0;
    SS1[12][3] = 4'h0;
    SS1[13][3] = 4'h0;
    SS1[14][3] = 4'h0;
    SS1[15][3] = 4'h0;
    SS1[16][3] = 4'hC;
    SS1[17][3] = 4'hC;
    SS1[18][3] = 4'hC;
    SS1[19][3] = 4'hC;
    SS1[20][3] = 4'hC;
    SS1[21][3] = 4'hD;
    SS1[22][3] = 4'hD;
    SS1[23][3] = 4'h0;
    SS1[24][3] = 4'h0;
    SS1[25][3] = 4'h0;
    SS1[26][3] = 4'h0;
    SS1[27][3] = 4'h0;
    SS1[28][3] = 4'h0;
    SS1[29][3] = 4'h0;
    SS1[30][3] = 4'h0;
    SS1[31][3] = 4'h0;
    SS1[32][3] = 4'h0;
    SS1[33][3] = 4'h0;
    SS1[34][3] = 4'h0;
    SS1[35][3] = 4'h0;
    SS1[36][3] = 4'h0;
    SS1[37][3] = 4'h0;
    SS1[38][3] = 4'h0;
    SS1[39][3] = 4'h0;
    SS1[40][3] = 4'h0;
    SS1[41][3] = 4'h0;
    SS1[42][3] = 4'h0;
    SS1[43][3] = 4'h0;
    SS1[44][3] = 4'h0;
    SS1[45][3] = 4'h0;
    SS1[46][3] = 4'h0;
    SS1[47][3] = 4'h0;
    SS1[0][4] = 4'h0;
    SS1[1][4] = 4'h0;
    SS1[2][4] = 4'h0;
    SS1[3][4] = 4'h0;
    SS1[4][4] = 4'h0;
    SS1[5][4] = 4'h0;
    SS1[6][4] = 4'h0;
    SS1[7][4] = 4'h0;
    SS1[8][4] = 4'h0;
    SS1[9][4] = 4'h0;
    SS1[10][4] = 4'h0;
    SS1[11][4] = 4'h0;
    SS1[12][4] = 4'h0;
    SS1[13][4] = 4'h0;
    SS1[14][4] = 4'h0;
    SS1[15][4] = 4'h0;
    SS1[16][4] = 4'hC;
    SS1[17][4] = 4'hC;
    SS1[18][4] = 4'hC;
    SS1[19][4] = 4'hC;
    SS1[20][4] = 4'hC;
    SS1[21][4] = 4'hC;
    SS1[22][4] = 4'hE;
    SS1[23][4] = 4'h0;
    SS1[24][4] = 4'h0;
    SS1[25][4] = 4'h0;
    SS1[26][4] = 4'h0;
    SS1[27][4] = 4'h0;
    SS1[28][4] = 4'h0;
    SS1[29][4] = 4'h0;
    SS1[30][4] = 4'h0;
    SS1[31][4] = 4'h0;
    SS1[32][4] = 4'h0;
    SS1[33][4] = 4'h0;
    SS1[34][4] = 4'h0;
    SS1[35][4] = 4'h0;
    SS1[36][4] = 4'h0;
    SS1[37][4] = 4'h0;
    SS1[38][4] = 4'h0;
    SS1[39][4] = 4'h0;
    SS1[40][4] = 4'h0;
    SS1[41][4] = 4'h0;
    SS1[42][4] = 4'h0;
    SS1[43][4] = 4'h0;
    SS1[44][4] = 4'h0;
    SS1[45][4] = 4'h0;
    SS1[46][4] = 4'h0;
    SS1[47][4] = 4'h0;
    SS1[0][5] = 4'h0;
    SS1[1][5] = 4'h0;
    SS1[2][5] = 4'h0;
    SS1[3][5] = 4'h0;
    SS1[4][5] = 4'h0;
    SS1[5][5] = 4'h0;
    SS1[6][5] = 4'h0;
    SS1[7][5] = 4'h0;
    SS1[8][5] = 4'h0;
    SS1[9][5] = 4'h0;
    SS1[10][5] = 4'h0;
    SS1[11][5] = 4'h0;
    SS1[12][5] = 4'h0;
    SS1[13][5] = 4'h0;
    SS1[14][5] = 4'h0;
    SS1[15][5] = 4'h0;
    SS1[16][5] = 4'h0;
    SS1[17][5] = 4'h0;
    SS1[18][5] = 4'hC;
    SS1[19][5] = 4'hC;
    SS1[20][5] = 4'hC;
    SS1[21][5] = 4'hC;
    SS1[22][5] = 4'hE;
    SS1[23][5] = 4'hE;
    SS1[24][5] = 4'hE;
    SS1[25][5] = 4'h0;
    SS1[26][5] = 4'h0;
    SS1[27][5] = 4'h0;
    SS1[28][5] = 4'h0;
    SS1[29][5] = 4'h0;
    SS1[30][5] = 4'h0;
    SS1[31][5] = 4'h0;
    SS1[32][5] = 4'h0;
    SS1[33][5] = 4'h0;
    SS1[34][5] = 4'h0;
    SS1[35][5] = 4'h0;
    SS1[36][5] = 4'h0;
    SS1[37][5] = 4'h0;
    SS1[38][5] = 4'h0;
    SS1[39][5] = 4'h0;
    SS1[40][5] = 4'h0;
    SS1[41][5] = 4'h0;
    SS1[42][5] = 4'h0;
    SS1[43][5] = 4'h0;
    SS1[44][5] = 4'h0;
    SS1[45][5] = 4'h0;
    SS1[46][5] = 4'h0;
    SS1[47][5] = 4'h0;
    SS1[0][6] = 4'h0;
    SS1[1][6] = 4'h0;
    SS1[2][6] = 4'h0;
    SS1[3][6] = 4'h0;
    SS1[4][6] = 4'h0;
    SS1[5][6] = 4'h0;
    SS1[6][6] = 4'h0;
    SS1[7][6] = 4'h0;
    SS1[8][6] = 4'h0;
    SS1[9][6] = 4'h0;
    SS1[10][6] = 4'h0;
    SS1[11][6] = 4'h0;
    SS1[12][6] = 4'h0;
    SS1[13][6] = 4'h0;
    SS1[14][6] = 4'h0;
    SS1[15][6] = 4'h0;
    SS1[16][6] = 4'h0;
    SS1[17][6] = 4'h0;
    SS1[18][6] = 4'hC;
    SS1[19][6] = 4'hC;
    SS1[20][6] = 4'hC;
    SS1[21][6] = 4'hC;
    SS1[22][6] = 4'hE;
    SS1[23][6] = 4'hE;
    SS1[24][6] = 4'hE;
    SS1[25][6] = 4'h0;
    SS1[26][6] = 4'h0;
    SS1[27][6] = 4'h0;
    SS1[28][6] = 4'h0;
    SS1[29][6] = 4'h0;
    SS1[30][6] = 4'h0;
    SS1[31][6] = 4'h0;
    SS1[32][6] = 4'h0;
    SS1[33][6] = 4'h0;
    SS1[34][6] = 4'h0;
    SS1[35][6] = 4'h0;
    SS1[36][6] = 4'h0;
    SS1[37][6] = 4'h0;
    SS1[38][6] = 4'h0;
    SS1[39][6] = 4'h0;
    SS1[40][6] = 4'h0;
    SS1[41][6] = 4'h0;
    SS1[42][6] = 4'h0;
    SS1[43][6] = 4'h0;
    SS1[44][6] = 4'h0;
    SS1[45][6] = 4'h0;
    SS1[46][6] = 4'h0;
    SS1[47][6] = 4'h0;
    SS1[0][7] = 4'h0;
    SS1[1][7] = 4'h0;
    SS1[2][7] = 4'h0;
    SS1[3][7] = 4'h0;
    SS1[4][7] = 4'h0;
    SS1[5][7] = 4'hD;
    SS1[6][7] = 4'hD;
    SS1[7][7] = 4'h0;
    SS1[8][7] = 4'h0;
    SS1[9][7] = 4'h0;
    SS1[10][7] = 4'h0;
    SS1[11][7] = 4'h0;
    SS1[12][7] = 4'h0;
    SS1[13][7] = 4'h0;
    SS1[14][7] = 4'h0;
    SS1[15][7] = 4'h0;
    SS1[16][7] = 4'h0;
    SS1[17][7] = 4'h0;
    SS1[18][7] = 4'hC;
    SS1[19][7] = 4'hC;
    SS1[20][7] = 4'hC;
    SS1[21][7] = 4'hD;
    SS1[22][7] = 4'hD;
    SS1[23][7] = 4'hE;
    SS1[24][7] = 4'h0;
    SS1[25][7] = 4'h0;
    SS1[26][7] = 4'h0;
    SS1[27][7] = 4'h0;
    SS1[28][7] = 4'h0;
    SS1[29][7] = 4'h0;
    SS1[30][7] = 4'h0;
    SS1[31][7] = 4'h0;
    SS1[32][7] = 4'h0;
    SS1[33][7] = 4'h0;
    SS1[34][7] = 4'h0;
    SS1[35][7] = 4'h0;
    SS1[36][7] = 4'h0;
    SS1[37][7] = 4'h0;
    SS1[38][7] = 4'h0;
    SS1[39][7] = 4'h0;
    SS1[40][7] = 4'h0;
    SS1[41][7] = 4'h0;
    SS1[42][7] = 4'h0;
    SS1[43][7] = 4'h0;
    SS1[44][7] = 4'hD;
    SS1[45][7] = 4'hD;
    SS1[46][7] = 4'h0;
    SS1[47][7] = 4'h0;
    SS1[0][8] = 4'h0;
    SS1[1][8] = 4'h0;
    SS1[2][8] = 4'h0;
    SS1[3][8] = 4'h0;
    SS1[4][8] = 4'h0;
    SS1[5][8] = 4'hD;
    SS1[6][8] = 4'hD;
    SS1[7][8] = 4'hD;
    SS1[8][8] = 4'hD;
    SS1[9][8] = 4'hD;
    SS1[10][8] = 4'h0;
    SS1[11][8] = 4'h0;
    SS1[12][8] = 4'h0;
    SS1[13][8] = 4'h0;
    SS1[14][8] = 4'h0;
    SS1[15][8] = 4'h0;
    SS1[16][8] = 4'h0;
    SS1[17][8] = 4'h0;
    SS1[18][8] = 4'hC;
    SS1[19][8] = 4'hC;
    SS1[20][8] = 4'hC;
    SS1[21][8] = 4'hD;
    SS1[22][8] = 4'hD;
    SS1[23][8] = 4'hD;
    SS1[24][8] = 4'hE;
    SS1[25][8] = 4'h0;
    SS1[26][8] = 4'h0;
    SS1[27][8] = 4'h0;
    SS1[28][8] = 4'h0;
    SS1[29][8] = 4'h0;
    SS1[30][8] = 4'h0;
    SS1[31][8] = 4'h0;
    SS1[32][8] = 4'h0;
    SS1[33][8] = 4'h0;
    SS1[34][8] = 4'h0;
    SS1[35][8] = 4'h0;
    SS1[36][8] = 4'h0;
    SS1[37][8] = 4'h0;
    SS1[38][8] = 4'h0;
    SS1[39][8] = 4'h0;
    SS1[40][8] = 4'hD;
    SS1[41][8] = 4'h0;
    SS1[42][8] = 4'h0;
    SS1[43][8] = 4'hD;
    SS1[44][8] = 4'hD;
    SS1[45][8] = 4'hD;
    SS1[46][8] = 4'h0;
    SS1[47][8] = 4'h0;
    SS1[0][9] = 4'h0;
    SS1[1][9] = 4'h0;
    SS1[2][9] = 4'h0;
    SS1[3][9] = 4'h0;
    SS1[4][9] = 4'hD;
    SS1[5][9] = 4'hD;
    SS1[6][9] = 4'hD;
    SS1[7][9] = 4'hD;
    SS1[8][9] = 4'hD;
    SS1[9][9] = 4'hD;
    SS1[10][9] = 4'hD;
    SS1[11][9] = 4'hE;
    SS1[12][9] = 4'h0;
    SS1[13][9] = 4'h0;
    SS1[14][9] = 4'h0;
    SS1[15][9] = 4'h0;
    SS1[16][9] = 4'h0;
    SS1[17][9] = 4'hC;
    SS1[18][9] = 4'hC;
    SS1[19][9] = 4'hC;
    SS1[20][9] = 4'hD;
    SS1[21][9] = 4'hD;
    SS1[22][9] = 4'hD;
    SS1[23][9] = 4'hD;
    SS1[24][9] = 4'hE;
    SS1[25][9] = 4'hE;
    SS1[26][9] = 4'hE;
    SS1[27][9] = 4'h0;
    SS1[28][9] = 4'h0;
    SS1[29][9] = 4'h0;
    SS1[30][9] = 4'h0;
    SS1[31][9] = 4'h0;
    SS1[32][9] = 4'h0;
    SS1[33][9] = 4'h0;
    SS1[34][9] = 4'h0;
    SS1[35][9] = 4'h0;
    SS1[36][9] = 4'h0;
    SS1[37][9] = 4'h0;
    SS1[38][9] = 4'h0;
    SS1[39][9] = 4'h0;
    SS1[40][9] = 4'hD;
    SS1[41][9] = 4'hD;
    SS1[42][9] = 4'hD;
    SS1[43][9] = 4'hD;
    SS1[44][9] = 4'hD;
    SS1[45][9] = 4'hD;
    SS1[46][9] = 4'h0;
    SS1[47][9] = 4'h0;
    SS1[0][10] = 4'h0;
    SS1[1][10] = 4'h0;
    SS1[2][10] = 4'h0;
    SS1[3][10] = 4'h0;
    SS1[4][10] = 4'h0;
    SS1[5][10] = 4'h0;
    SS1[6][10] = 4'h0;
    SS1[7][10] = 4'hD;
    SS1[8][10] = 4'hD;
    SS1[9][10] = 4'hD;
    SS1[10][10] = 4'hE;
    SS1[11][10] = 4'hE;
    SS1[12][10] = 4'hE;
    SS1[13][10] = 4'hE;
    SS1[14][10] = 4'hE;
    SS1[15][10] = 4'h0;
    SS1[16][10] = 4'h0;
    SS1[17][10] = 4'hC;
    SS1[18][10] = 4'hC;
    SS1[19][10] = 4'hC;
    SS1[20][10] = 4'hC;
    SS1[21][10] = 4'hC;
    SS1[22][10] = 4'hD;
    SS1[23][10] = 4'hE;
    SS1[24][10] = 4'hE;
    SS1[25][10] = 4'hE;
    SS1[26][10] = 4'h0;
    SS1[27][10] = 4'h0;
    SS1[28][10] = 4'h0;
    SS1[29][10] = 4'h0;
    SS1[30][10] = 4'h0;
    SS1[31][10] = 4'h0;
    SS1[32][10] = 4'h0;
    SS1[33][10] = 4'h0;
    SS1[34][10] = 4'h0;
    SS1[35][10] = 4'h0;
    SS1[36][10] = 4'hE;
    SS1[37][10] = 4'hE;
    SS1[38][10] = 4'h0;
    SS1[39][10] = 4'hD;
    SS1[40][10] = 4'hD;
    SS1[41][10] = 4'hD;
    SS1[42][10] = 4'hC;
    SS1[43][10] = 4'hC;
    SS1[44][10] = 4'hC;
    SS1[45][10] = 4'hC;
    SS1[46][10] = 4'h0;
    SS1[47][10] = 4'h0;
    SS1[0][11] = 4'h0;
    SS1[1][11] = 4'h0;
    SS1[2][11] = 4'h0;
    SS1[3][11] = 4'h0;
    SS1[4][11] = 4'h0;
    SS1[5][11] = 4'h0;
    SS1[6][11] = 4'h0;
    SS1[7][11] = 4'hD;
    SS1[8][11] = 4'hD;
    SS1[9][11] = 4'hD;
    SS1[10][11] = 4'hE;
    SS1[11][11] = 4'hE;
    SS1[12][11] = 4'hE;
    SS1[13][11] = 4'hE;
    SS1[14][11] = 4'hE;
    SS1[15][11] = 4'hE;
    SS1[16][11] = 4'hC;
    SS1[17][11] = 4'hC;
    SS1[18][11] = 4'hC;
    SS1[19][11] = 4'hC;
    SS1[20][11] = 4'hC;
    SS1[21][11] = 4'hC;
    SS1[22][11] = 4'hC;
    SS1[23][11] = 4'hD;
    SS1[24][11] = 4'hD;
    SS1[25][11] = 4'hE;
    SS1[26][11] = 4'h0;
    SS1[27][11] = 4'h0;
    SS1[28][11] = 4'h0;
    SS1[29][11] = 4'h0;
    SS1[30][11] = 4'h0;
    SS1[31][11] = 4'h0;
    SS1[32][11] = 4'hE;
    SS1[33][11] = 4'h0;
    SS1[34][11] = 4'h0;
    SS1[35][11] = 4'h0;
    SS1[36][11] = 4'hE;
    SS1[37][11] = 4'hE;
    SS1[38][11] = 4'hE;
    SS1[39][11] = 4'hC;
    SS1[40][11] = 4'hD;
    SS1[41][11] = 4'hD;
    SS1[42][11] = 4'hC;
    SS1[43][11] = 4'hC;
    SS1[44][11] = 4'hC;
    SS1[45][11] = 4'h0;
    SS1[46][11] = 4'h0;
    SS1[47][11] = 4'h0;
    SS1[0][12] = 4'h0;
    SS1[1][12] = 4'h0;
    SS1[2][12] = 4'h0;
    SS1[3][12] = 4'h0;
    SS1[4][12] = 4'h0;
    SS1[5][12] = 4'h0;
    SS1[6][12] = 4'hD;
    SS1[7][12] = 4'hD;
    SS1[8][12] = 4'hD;
    SS1[9][12] = 4'hD;
    SS1[10][12] = 4'hD;
    SS1[11][12] = 4'hD;
    SS1[12][12] = 4'hE;
    SS1[13][12] = 4'hE;
    SS1[14][12] = 4'hE;
    SS1[15][12] = 4'hE;
    SS1[16][12] = 4'hC;
    SS1[17][12] = 4'hC;
    SS1[18][12] = 4'hC;
    SS1[19][12] = 4'hC;
    SS1[20][12] = 4'hC;
    SS1[21][12] = 4'hC;
    SS1[22][12] = 4'hD;
    SS1[23][12] = 4'hD;
    SS1[24][12] = 4'hD;
    SS1[25][12] = 4'hD;
    SS1[26][12] = 4'hE;
    SS1[27][12] = 4'h0;
    SS1[28][12] = 4'h0;
    SS1[29][12] = 4'h0;
    SS1[30][12] = 4'h0;
    SS1[31][12] = 4'h0;
    SS1[32][12] = 4'hE;
    SS1[33][12] = 4'hE;
    SS1[34][12] = 4'hE;
    SS1[35][12] = 4'hE;
    SS1[36][12] = 4'hE;
    SS1[37][12] = 4'hE;
    SS1[38][12] = 4'hC;
    SS1[39][12] = 4'hC;
    SS1[40][12] = 4'hC;
    SS1[41][12] = 4'hC;
    SS1[42][12] = 4'hC;
    SS1[43][12] = 4'hC;
    SS1[44][12] = 4'hC;
    SS1[45][12] = 4'h0;
    SS1[46][12] = 4'h0;
    SS1[47][12] = 4'h0;
    SS1[0][13] = 4'h0;
    SS1[1][13] = 4'h0;
    SS1[2][13] = 4'h0;
    SS1[3][13] = 4'h0;
    SS1[4][13] = 4'h0;
    SS1[5][13] = 4'h0;
    SS1[6][13] = 4'hD;
    SS1[7][13] = 4'hD;
    SS1[8][13] = 4'hD;
    SS1[9][13] = 4'hD;
    SS1[10][13] = 4'hD;
    SS1[11][13] = 4'hD;
    SS1[12][13] = 4'hE;
    SS1[13][13] = 4'hE;
    SS1[14][13] = 4'hE;
    SS1[15][13] = 4'hE;
    SS1[16][13] = 4'hC;
    SS1[17][13] = 4'hC;
    SS1[18][13] = 4'hC;
    SS1[19][13] = 4'hC;
    SS1[20][13] = 4'hC;
    SS1[21][13] = 4'hC;
    SS1[22][13] = 4'hD;
    SS1[23][13] = 4'hD;
    SS1[24][13] = 4'hD;
    SS1[25][13] = 4'hE;
    SS1[26][13] = 4'hE;
    SS1[27][13] = 4'hE;
    SS1[28][13] = 4'hE;
    SS1[29][13] = 4'hE;
    SS1[30][13] = 4'h0;
    SS1[31][13] = 4'h0;
    SS1[32][13] = 4'hE;
    SS1[33][13] = 4'hE;
    SS1[34][13] = 4'hE;
    SS1[35][13] = 4'hD;
    SS1[36][13] = 4'hD;
    SS1[37][13] = 4'hE;
    SS1[38][13] = 4'hC;
    SS1[39][13] = 4'hC;
    SS1[40][13] = 4'hC;
    SS1[41][13] = 4'hC;
    SS1[42][13] = 4'hC;
    SS1[43][13] = 4'hC;
    SS1[44][13] = 4'h0;
    SS1[45][13] = 4'h0;
    SS1[46][13] = 4'h0;
    SS1[47][13] = 4'h0;
    SS1[0][14] = 4'h0;
    SS1[1][14] = 4'h0;
    SS1[2][14] = 4'h0;
    SS1[3][14] = 4'h0;
    SS1[4][14] = 4'h0;
    SS1[5][14] = 4'h0;
    SS1[6][14] = 4'h0;
    SS1[7][14] = 4'h0;
    SS1[8][14] = 4'h0;
    SS1[9][14] = 4'hD;
    SS1[10][14] = 4'hD;
    SS1[11][14] = 4'hD;
    SS1[12][14] = 4'hE;
    SS1[13][14] = 4'hE;
    SS1[14][14] = 4'hE;
    SS1[15][14] = 4'hE;
    SS1[16][14] = 4'hE;
    SS1[17][14] = 4'hC;
    SS1[18][14] = 4'hC;
    SS1[19][14] = 4'hC;
    SS1[20][14] = 4'hC;
    SS1[21][14] = 4'hC;
    SS1[22][14] = 4'hC;
    SS1[23][14] = 4'hC;
    SS1[24][14] = 4'hD;
    SS1[25][14] = 4'hE;
    SS1[26][14] = 4'hE;
    SS1[27][14] = 4'hE;
    SS1[28][14] = 4'hE;
    SS1[29][14] = 4'hE;
    SS1[30][14] = 4'hE;
    SS1[31][14] = 4'hD;
    SS1[32][14] = 4'hE;
    SS1[33][14] = 4'hE;
    SS1[34][14] = 4'hD;
    SS1[35][14] = 4'hD;
    SS1[36][14] = 4'hD;
    SS1[37][14] = 4'hD;
    SS1[38][14] = 4'hC;
    SS1[39][14] = 4'hC;
    SS1[40][14] = 4'hC;
    SS1[41][14] = 4'hC;
    SS1[42][14] = 4'hC;
    SS1[43][14] = 4'hC;
    SS1[44][14] = 4'h0;
    SS1[45][14] = 4'h0;
    SS1[46][14] = 4'h0;
    SS1[47][14] = 4'h0;
    SS1[0][15] = 4'h0;
    SS1[1][15] = 4'h0;
    SS1[2][15] = 4'h0;
    SS1[3][15] = 4'h0;
    SS1[4][15] = 4'h0;
    SS1[5][15] = 4'h0;
    SS1[6][15] = 4'h0;
    SS1[7][15] = 4'h0;
    SS1[8][15] = 4'h3;
    SS1[9][15] = 4'h3;
    SS1[10][15] = 4'h3;
    SS1[11][15] = 4'hE;
    SS1[12][15] = 4'hE;
    SS1[13][15] = 4'hE;
    SS1[14][15] = 4'hE;
    SS1[15][15] = 4'hE;
    SS1[16][15] = 4'hE;
    SS1[17][15] = 4'hE;
    SS1[18][15] = 4'hC;
    SS1[19][15] = 4'hC;
    SS1[20][15] = 4'hC;
    SS1[21][15] = 4'hC;
    SS1[22][15] = 4'hC;
    SS1[23][15] = 4'hC;
    SS1[24][15] = 4'hE;
    SS1[25][15] = 4'hE;
    SS1[26][15] = 4'hE;
    SS1[27][15] = 4'hE;
    SS1[28][15] = 4'hE;
    SS1[29][15] = 4'hE;
    SS1[30][15] = 4'hE;
    SS1[31][15] = 4'hD;
    SS1[32][15] = 4'hD;
    SS1[33][15] = 4'hD;
    SS1[34][15] = 4'hD;
    SS1[35][15] = 4'hD;
    SS1[36][15] = 4'hD;
    SS1[37][15] = 4'hC;
    SS1[38][15] = 4'hC;
    SS1[39][15] = 4'hC;
    SS1[40][15] = 4'h0;
    SS1[41][15] = 4'h0;
    SS1[42][15] = 4'hC;
    SS1[43][15] = 4'hC;
    SS1[44][15] = 4'h0;
    SS1[45][15] = 4'h0;
    SS1[46][15] = 4'h0;
    SS1[47][15] = 4'h0;
    SS1[0][16] = 4'h0;
    SS1[1][16] = 4'h0;
    SS1[2][16] = 4'h0;
    SS1[3][16] = 4'h0;
    SS1[4][16] = 4'h0;
    SS1[5][16] = 4'h0;
    SS1[6][16] = 4'h0;
    SS1[7][16] = 4'h0;
    SS1[8][16] = 4'h3;
    SS1[9][16] = 4'h3;
    SS1[10][16] = 4'h3;
    SS1[11][16] = 4'hD;
    SS1[12][16] = 4'hD;
    SS1[13][16] = 4'hD;
    SS1[14][16] = 4'hE;
    SS1[15][16] = 4'hE;
    SS1[16][16] = 4'hE;
    SS1[17][16] = 4'hC;
    SS1[18][16] = 4'hC;
    SS1[19][16] = 4'hC;
    SS1[20][16] = 4'hC;
    SS1[21][16] = 4'hC;
    SS1[22][16] = 4'hC;
    SS1[23][16] = 4'hC;
    SS1[24][16] = 4'hE;
    SS1[25][16] = 4'hE;
    SS1[26][16] = 4'hE;
    SS1[27][16] = 4'hE;
    SS1[28][16] = 4'hE;
    SS1[29][16] = 4'hE;
    SS1[30][16] = 4'hD;
    SS1[31][16] = 4'hD;
    SS1[32][16] = 4'hD;
    SS1[33][16] = 4'hD;
    SS1[34][16] = 4'hC;
    SS1[35][16] = 4'hC;
    SS1[36][16] = 4'hC;
    SS1[37][16] = 4'hC;
    SS1[38][16] = 4'hC;
    SS1[39][16] = 4'hC;
    SS1[40][16] = 4'h0;
    SS1[41][16] = 4'h0;
    SS1[42][16] = 4'h0;
    SS1[43][16] = 4'h0;
    SS1[44][16] = 4'h0;
    SS1[45][16] = 4'h0;
    SS1[46][16] = 4'h0;
    SS1[47][16] = 4'h0;
    SS1[0][17] = 4'h0;
    SS1[1][17] = 4'h0;
    SS1[2][17] = 4'h0;
    SS1[3][17] = 4'h0;
    SS1[4][17] = 4'h0;
    SS1[5][17] = 4'h0;
    SS1[6][17] = 4'h0;
    SS1[7][17] = 4'h0;
    SS1[8][17] = 4'h3;
    SS1[9][17] = 4'h3;
    SS1[10][17] = 4'h3;
    SS1[11][17] = 4'hD;
    SS1[12][17] = 4'hD;
    SS1[13][17] = 4'hD;
    SS1[14][17] = 4'hD;
    SS1[15][17] = 4'hD;
    SS1[16][17] = 4'hE;
    SS1[17][17] = 4'hC;
    SS1[18][17] = 4'hC;
    SS1[19][17] = 4'hC;
    SS1[20][17] = 4'hC;
    SS1[21][17] = 4'hC;
    SS1[22][17] = 4'hC;
    SS1[23][17] = 4'hD;
    SS1[24][17] = 4'hE;
    SS1[25][17] = 4'hE;
    SS1[26][17] = 4'hE;
    SS1[27][17] = 4'hE;
    SS1[28][17] = 4'hE;
    SS1[29][17] = 4'hE;
    SS1[30][17] = 4'hC;
    SS1[31][17] = 4'hC;
    SS1[32][17] = 4'hD;
    SS1[33][17] = 4'hC;
    SS1[34][17] = 4'hC;
    SS1[35][17] = 4'hC;
    SS1[36][17] = 4'hC;
    SS1[37][17] = 4'hC;
    SS1[38][17] = 4'hC;
    SS1[39][17] = 4'hC;
    SS1[40][17] = 4'h0;
    SS1[41][17] = 4'h0;
    SS1[42][17] = 4'h0;
    SS1[43][17] = 4'h0;
    SS1[44][17] = 4'h0;
    SS1[45][17] = 4'h0;
    SS1[46][17] = 4'h0;
    SS1[47][17] = 4'h0;
    SS1[0][18] = 4'h0;
    SS1[1][18] = 4'h0;
    SS1[2][18] = 4'h0;
    SS1[3][18] = 4'h0;
    SS1[4][18] = 4'h0;
    SS1[5][18] = 4'h0;
    SS1[6][18] = 4'h0;
    SS1[7][18] = 4'h0;
    SS1[8][18] = 4'h0;
    SS1[9][18] = 4'h0;
    SS1[10][18] = 4'h0;
    SS1[11][18] = 4'hD;
    SS1[12][18] = 4'hD;
    SS1[13][18] = 4'hD;
    SS1[14][18] = 4'hD;
    SS1[15][18] = 4'hD;
    SS1[16][18] = 4'hD;
    SS1[17][18] = 4'hE;
    SS1[18][18] = 4'hC;
    SS1[19][18] = 4'hC;
    SS1[20][18] = 4'hC;
    SS1[21][18] = 4'hC;
    SS1[22][18] = 4'hC;
    SS1[23][18] = 4'hD;
    SS1[24][18] = 4'hD;
    SS1[25][18] = 4'hD;
    SS1[26][18] = 4'hE;
    SS1[27][18] = 4'hE;
    SS1[28][18] = 4'hE;
    SS1[29][18] = 4'hC;
    SS1[30][18] = 4'hC;
    SS1[31][18] = 4'hC;
    SS1[32][18] = 4'hC;
    SS1[33][18] = 4'hC;
    SS1[34][18] = 4'hC;
    SS1[35][18] = 4'hC;
    SS1[36][18] = 4'hC;
    SS1[37][18] = 4'hC;
    SS1[38][18] = 4'hC;
    SS1[39][18] = 4'h0;
    SS1[40][18] = 4'h0;
    SS1[41][18] = 4'h0;
    SS1[42][18] = 4'h0;
    SS1[43][18] = 4'h0;
    SS1[44][18] = 4'h0;
    SS1[45][18] = 4'h0;
    SS1[46][18] = 4'h0;
    SS1[47][18] = 4'h0;
    SS1[0][19] = 4'h0;
    SS1[1][19] = 4'h0;
    SS1[2][19] = 4'h0;
    SS1[3][19] = 4'h0;
    SS1[4][19] = 4'h0;
    SS1[5][19] = 4'h0;
    SS1[6][19] = 4'h0;
    SS1[7][19] = 4'h0;
    SS1[8][19] = 4'h0;
    SS1[9][19] = 4'h0;
    SS1[10][19] = 4'h0;
    SS1[11][19] = 4'h0;
    SS1[12][19] = 4'h0;
    SS1[13][19] = 4'hD;
    SS1[14][19] = 4'hD;
    SS1[15][19] = 4'hD;
    SS1[16][19] = 4'hE;
    SS1[17][19] = 4'hE;
    SS1[18][19] = 4'hE;
    SS1[19][19] = 4'hC;
    SS1[20][19] = 4'hC;
    SS1[21][19] = 4'hC;
    SS1[22][19] = 4'hC;
    SS1[23][19] = 4'hD;
    SS1[24][19] = 4'hD;
    SS1[25][19] = 4'hD;
    SS1[26][19] = 4'hD;
    SS1[27][19] = 4'hD;
    SS1[28][19] = 4'hD;
    SS1[29][19] = 4'hC;
    SS1[30][19] = 4'hC;
    SS1[31][19] = 4'hC;
    SS1[32][19] = 4'hC;
    SS1[33][19] = 4'hC;
    SS1[34][19] = 4'hC;
    SS1[35][19] = 4'hC;
    SS1[36][19] = 4'hC;
    SS1[37][19] = 4'hC;
    SS1[38][19] = 4'hC;
    SS1[39][19] = 4'h0;
    SS1[40][19] = 4'h0;
    SS1[41][19] = 4'h0;
    SS1[42][19] = 4'h0;
    SS1[43][19] = 4'h0;
    SS1[44][19] = 4'h0;
    SS1[45][19] = 4'h0;
    SS1[46][19] = 4'h0;
    SS1[47][19] = 4'h0;
    SS1[0][20] = 4'h0;
    SS1[1][20] = 4'h0;
    SS1[2][20] = 4'h0;
    SS1[3][20] = 4'h0;
    SS1[4][20] = 4'h0;
    SS1[5][20] = 4'h0;
    SS1[6][20] = 4'h0;
    SS1[7][20] = 4'h0;
    SS1[8][20] = 4'h0;
    SS1[9][20] = 4'h0;
    SS1[10][20] = 4'h0;
    SS1[11][20] = 4'h0;
    SS1[12][20] = 4'h0;
    SS1[13][20] = 4'hD;
    SS1[14][20] = 4'hD;
    SS1[15][20] = 4'hD;
    SS1[16][20] = 4'hE;
    SS1[17][20] = 4'hE;
    SS1[18][20] = 4'hE;
    SS1[19][20] = 4'hC;
    SS1[20][20] = 4'hC;
    SS1[21][20] = 4'hC;
    SS1[22][20] = 4'hC;
    SS1[23][20] = 4'hD;
    SS1[24][20] = 4'hD;
    SS1[25][20] = 4'hD;
    SS1[26][20] = 4'hD;
    SS1[27][20] = 4'hD;
    SS1[28][20] = 4'hD;
    SS1[29][20] = 4'hC;
    SS1[30][20] = 4'hC;
    SS1[31][20] = 4'hC;
    SS1[32][20] = 4'hC;
    SS1[33][20] = 4'hC;
    SS1[34][20] = 4'hC;
    SS1[35][20] = 4'hC;
    SS1[36][20] = 4'hC;
    SS1[37][20] = 4'hC;
    SS1[38][20] = 4'hE;
    SS1[39][20] = 4'h0;
    SS1[40][20] = 4'h0;
    SS1[41][20] = 4'h0;
    SS1[42][20] = 4'h0;
    SS1[43][20] = 4'h0;
    SS1[44][20] = 4'h0;
    SS1[45][20] = 4'h0;
    SS1[46][20] = 4'h0;
    SS1[47][20] = 4'h0;
    SS1[0][21] = 4'h0;
    SS1[1][21] = 4'h0;
    SS1[2][21] = 4'h0;
    SS1[3][21] = 4'h0;
    SS1[4][21] = 4'h0;
    SS1[5][21] = 4'h0;
    SS1[6][21] = 4'h0;
    SS1[7][21] = 4'h0;
    SS1[8][21] = 4'h0;
    SS1[9][21] = 4'h0;
    SS1[10][21] = 4'h0;
    SS1[11][21] = 4'h0;
    SS1[12][21] = 4'hD;
    SS1[13][21] = 4'hD;
    SS1[14][21] = 4'hD;
    SS1[15][21] = 4'hD;
    SS1[16][21] = 4'hD;
    SS1[17][21] = 4'hD;
    SS1[18][21] = 4'hE;
    SS1[19][21] = 4'hC;
    SS1[20][21] = 4'hC;
    SS1[21][21] = 4'hC;
    SS1[22][21] = 4'hC;
    SS1[23][21] = 4'hC;
    SS1[24][21] = 4'hC;
    SS1[25][21] = 4'hC;
    SS1[26][21] = 4'hD;
    SS1[27][21] = 4'hD;
    SS1[28][21] = 4'hC;
    SS1[29][21] = 4'hC;
    SS1[30][21] = 4'hC;
    SS1[31][21] = 4'hC;
    SS1[32][21] = 4'hC;
    SS1[33][21] = 4'hC;
    SS1[34][21] = 4'hC;
    SS1[35][21] = 4'hC;
    SS1[36][21] = 4'hC;
    SS1[37][21] = 4'hC;
    SS1[38][21] = 4'hE;
    SS1[39][21] = 4'hE;
    SS1[40][21] = 4'hE;
    SS1[41][21] = 4'h0;
    SS1[42][21] = 4'h0;
    SS1[43][21] = 4'h0;
    SS1[44][21] = 4'h0;
    SS1[45][21] = 4'h0;
    SS1[46][21] = 4'h0;
    SS1[47][21] = 4'h0;
    SS1[0][22] = 4'h0;
    SS1[1][22] = 4'h0;
    SS1[2][22] = 4'h0;
    SS1[3][22] = 4'h0;
    SS1[4][22] = 4'h0;
    SS1[5][22] = 4'h0;
    SS1[6][22] = 4'h0;
    SS1[7][22] = 4'h0;
    SS1[8][22] = 4'h0;
    SS1[9][22] = 4'h0;
    SS1[10][22] = 4'h0;
    SS1[11][22] = 4'h0;
    SS1[12][22] = 4'h3;
    SS1[13][22] = 4'hD;
    SS1[14][22] = 4'hD;
    SS1[15][22] = 4'hD;
    SS1[16][22] = 4'hD;
    SS1[17][22] = 4'hD;
    SS1[18][22] = 4'hC;
    SS1[19][22] = 4'hC;
    SS1[20][22] = 4'hC;
    SS1[21][22] = 4'hC;
    SS1[22][22] = 4'hC;
    SS1[23][22] = 4'hC;
    SS1[24][22] = 4'hC;
    SS1[25][22] = 4'hC;
    SS1[26][22] = 4'hC;
    SS1[27][22] = 4'hC;
    SS1[28][22] = 4'hC;
    SS1[29][22] = 4'hC;
    SS1[30][22] = 4'hC;
    SS1[31][22] = 4'hC;
    SS1[32][22] = 4'hC;
    SS1[33][22] = 4'hC;
    SS1[34][22] = 4'hE;
    SS1[35][22] = 4'hE;
    SS1[36][22] = 4'hC;
    SS1[37][22] = 4'hE;
    SS1[38][22] = 4'hE;
    SS1[39][22] = 4'hE;
    SS1[40][22] = 4'hE;
    SS1[41][22] = 4'hE;
    SS1[42][22] = 4'hE;
    SS1[43][22] = 4'hE;
    SS1[44][22] = 4'h0;
    SS1[45][22] = 4'h0;
    SS1[46][22] = 4'h0;
    SS1[47][22] = 4'h0;
    SS1[0][23] = 4'h0;
    SS1[1][23] = 4'h0;
    SS1[2][23] = 4'h0;
    SS1[3][23] = 4'h0;
    SS1[4][23] = 4'h0;
    SS1[5][23] = 4'h0;
    SS1[6][23] = 4'h0;
    SS1[7][23] = 4'h0;
    SS1[8][23] = 4'h0;
    SS1[9][23] = 4'h0;
    SS1[10][23] = 4'h0;
    SS1[11][23] = 4'h3;
    SS1[12][23] = 4'h3;
    SS1[13][23] = 4'h3;
    SS1[14][23] = 4'h3;
    SS1[15][23] = 4'hD;
    SS1[16][23] = 4'hD;
    SS1[17][23] = 4'hD;
    SS1[18][23] = 4'hC;
    SS1[19][23] = 4'hC;
    SS1[20][23] = 4'hC;
    SS1[21][23] = 4'hD;
    SS1[22][23] = 4'hD;
    SS1[23][23] = 4'hC;
    SS1[24][23] = 4'hC;
    SS1[25][23] = 4'hC;
    SS1[26][23] = 4'hC;
    SS1[27][23] = 4'hC;
    SS1[28][23] = 4'hC;
    SS1[29][23] = 4'hC;
    SS1[30][23] = 4'hC;
    SS1[31][23] = 4'hC;
    SS1[32][23] = 4'hC;
    SS1[33][23] = 4'hC;
    SS1[34][23] = 4'hE;
    SS1[35][23] = 4'hE;
    SS1[36][23] = 4'hE;
    SS1[37][23] = 4'hE;
    SS1[38][23] = 4'hE;
    SS1[39][23] = 4'hE;
    SS1[40][23] = 4'hE;
    SS1[41][23] = 4'hE;
    SS1[42][23] = 4'hE;
    SS1[43][23] = 4'hD;
    SS1[44][23] = 4'hD;
    SS1[45][23] = 4'hD;
    SS1[46][23] = 4'h0;
    SS1[47][23] = 4'h0;
    SS1[0][24] = 4'h0;
    SS1[1][24] = 4'h0;
    SS1[2][24] = 4'h0;
    SS1[3][24] = 4'h0;
    SS1[4][24] = 4'h0;
    SS1[5][24] = 4'h0;
    SS1[6][24] = 4'h0;
    SS1[7][24] = 4'h0;
    SS1[8][24] = 4'h0;
    SS1[9][24] = 4'h0;
    SS1[10][24] = 4'h0;
    SS1[11][24] = 4'h3;
    SS1[12][24] = 4'h3;
    SS1[13][24] = 4'h3;
    SS1[14][24] = 4'hD;
    SS1[15][24] = 4'hD;
    SS1[16][24] = 4'hD;
    SS1[17][24] = 4'hC;
    SS1[18][24] = 4'hC;
    SS1[19][24] = 4'hC;
    SS1[20][24] = 4'hC;
    SS1[21][24] = 4'hD;
    SS1[22][24] = 4'hD;
    SS1[23][24] = 4'hD;
    SS1[24][24] = 4'hD;
    SS1[25][24] = 4'hC;
    SS1[26][24] = 4'hC;
    SS1[27][24] = 4'hC;
    SS1[28][24] = 4'hC;
    SS1[29][24] = 4'hC;
    SS1[30][24] = 4'hE;
    SS1[31][24] = 4'hE;
    SS1[32][24] = 4'hE;
    SS1[33][24] = 4'hE;
    SS1[34][24] = 4'hE;
    SS1[35][24] = 4'hE;
    SS1[36][24] = 4'hE;
    SS1[37][24] = 4'hE;
    SS1[38][24] = 4'hE;
    SS1[39][24] = 4'hE;
    SS1[40][24] = 4'hD;
    SS1[41][24] = 4'hE;
    SS1[42][24] = 4'hE;
    SS1[43][24] = 4'hD;
    SS1[44][24] = 4'hD;
    SS1[45][24] = 4'hD;
    SS1[46][24] = 4'hD;
    SS1[47][24] = 4'hD;
    SS1[0][25] = 4'h0;
    SS1[1][25] = 4'h0;
    SS1[2][25] = 4'h0;
    SS1[3][25] = 4'h0;
    SS1[4][25] = 4'h0;
    SS1[5][25] = 4'h0;
    SS1[6][25] = 4'h0;
    SS1[7][25] = 4'h0;
    SS1[8][25] = 4'h0;
    SS1[9][25] = 4'h0;
    SS1[10][25] = 4'h0;
    SS1[11][25] = 4'h0;
    SS1[12][25] = 4'h3;
    SS1[13][25] = 4'h3;
    SS1[14][25] = 4'hD;
    SS1[15][25] = 4'hD;
    SS1[16][25] = 4'hD;
    SS1[17][25] = 4'hD;
    SS1[18][25] = 4'hD;
    SS1[19][25] = 4'hD;
    SS1[20][25] = 4'hD;
    SS1[21][25] = 4'hD;
    SS1[22][25] = 4'hD;
    SS1[23][25] = 4'hD;
    SS1[24][25] = 4'hD;
    SS1[25][25] = 4'hD;
    SS1[26][25] = 4'hD;
    SS1[27][25] = 4'hC;
    SS1[28][25] = 4'hC;
    SS1[29][25] = 4'hC;
    SS1[30][25] = 4'hE;
    SS1[31][25] = 4'hE;
    SS1[32][25] = 4'hE;
    SS1[33][25] = 4'hD;
    SS1[34][25] = 4'hD;
    SS1[35][25] = 4'hE;
    SS1[36][25] = 4'hE;
    SS1[37][25] = 4'hE;
    SS1[38][25] = 4'hE;
    SS1[39][25] = 4'hD;
    SS1[40][25] = 4'hD;
    SS1[41][25] = 4'hD;
    SS1[42][25] = 4'hD;
    SS1[43][25] = 4'hD;
    SS1[44][25] = 4'hD;
    SS1[45][25] = 4'hD;
    SS1[46][25] = 4'hD;
    SS1[47][25] = 4'hD;
    SS1[0][26] = 4'h0;
    SS1[1][26] = 4'h0;
    SS1[2][26] = 4'h0;
    SS1[3][26] = 4'h0;
    SS1[4][26] = 4'h0;
    SS1[5][26] = 4'h0;
    SS1[6][26] = 4'h0;
    SS1[7][26] = 4'h0;
    SS1[8][26] = 4'h0;
    SS1[9][26] = 4'h0;
    SS1[10][26] = 4'h0;
    SS1[11][26] = 4'h0;
    SS1[12][26] = 4'h0;
    SS1[13][26] = 4'h0;
    SS1[14][26] = 4'hF;
    SS1[15][26] = 4'hD;
    SS1[16][26] = 4'hD;
    SS1[17][26] = 4'hD;
    SS1[18][26] = 4'hD;
    SS1[19][26] = 4'hD;
    SS1[20][26] = 4'hA;
    SS1[21][26] = 4'hA;
    SS1[22][26] = 4'hD;
    SS1[23][26] = 4'hD;
    SS1[24][26] = 4'hD;
    SS1[25][26] = 4'hD;
    SS1[26][26] = 4'hC;
    SS1[27][26] = 4'hC;
    SS1[28][26] = 4'hC;
    SS1[29][26] = 4'hD;
    SS1[30][26] = 4'hE;
    SS1[31][26] = 4'hE;
    SS1[32][26] = 4'hE;
    SS1[33][26] = 4'hD;
    SS1[34][26] = 4'hD;
    SS1[35][26] = 4'hD;
    SS1[36][26] = 4'hD;
    SS1[37][26] = 4'hD;
    SS1[38][26] = 4'hE;
    SS1[39][26] = 4'hD;
    SS1[40][26] = 4'hD;
    SS1[41][26] = 4'hD;
    SS1[42][26] = 4'hD;
    SS1[43][26] = 4'hD;
    SS1[44][26] = 4'hD;
    SS1[45][26] = 4'hE;
    SS1[46][26] = 4'hD;
    SS1[47][26] = 4'hD;
    SS1[0][27] = 4'h0;
    SS1[1][27] = 4'h0;
    SS1[2][27] = 4'h0;
    SS1[3][27] = 4'h0;
    SS1[4][27] = 4'h0;
    SS1[5][27] = 4'h0;
    SS1[6][27] = 4'h0;
    SS1[7][27] = 4'h0;
    SS1[8][27] = 4'h0;
    SS1[9][27] = 4'h0;
    SS1[10][27] = 4'h0;
    SS1[11][27] = 4'h0;
    SS1[12][27] = 4'h0;
    SS1[13][27] = 4'h0;
    SS1[14][27] = 4'h0;
    SS1[15][27] = 4'h0;
    SS1[16][27] = 4'hC;
    SS1[17][27] = 4'hD;
    SS1[18][27] = 4'hD;
    SS1[19][27] = 4'hA;
    SS1[20][27] = 4'hA;
    SS1[21][27] = 4'hA;
    SS1[22][27] = 4'hA;
    SS1[23][27] = 4'hA;
    SS1[24][27] = 4'hA;
    SS1[25][27] = 4'hD;
    SS1[26][27] = 4'hC;
    SS1[27][27] = 4'hC;
    SS1[28][27] = 4'hC;
    SS1[29][27] = 4'hD;
    SS1[30][27] = 4'hD;
    SS1[31][27] = 4'hD;
    SS1[32][27] = 4'hD;
    SS1[33][27] = 4'hD;
    SS1[34][27] = 4'hD;
    SS1[35][27] = 4'hD;
    SS1[36][27] = 4'hD;
    SS1[37][27] = 4'hD;
    SS1[38][27] = 4'hD;
    SS1[39][27] = 4'h3;
    SS1[40][27] = 4'hD;
    SS1[41][27] = 4'hD;
    SS1[42][27] = 4'hD;
    SS1[43][27] = 4'hD;
    SS1[44][27] = 4'hD;
    SS1[45][27] = 4'h0;
    SS1[46][27] = 4'h0;
    SS1[47][27] = 4'h0;
    SS1[0][28] = 4'h0;
    SS1[1][28] = 4'h0;
    SS1[2][28] = 4'h0;
    SS1[3][28] = 4'h0;
    SS1[4][28] = 4'h0;
    SS1[5][28] = 4'h0;
    SS1[6][28] = 4'h0;
    SS1[7][28] = 4'h0;
    SS1[8][28] = 4'h0;
    SS1[9][28] = 4'h0;
    SS1[10][28] = 4'h0;
    SS1[11][28] = 4'h0;
    SS1[12][28] = 4'h0;
    SS1[13][28] = 4'h0;
    SS1[14][28] = 4'h0;
    SS1[15][28] = 4'h0;
    SS1[16][28] = 4'hC;
    SS1[17][28] = 4'hC;
    SS1[18][28] = 4'hC;
    SS1[19][28] = 4'hA;
    SS1[20][28] = 4'hA;
    SS1[21][28] = 4'hA;
    SS1[22][28] = 4'hA;
    SS1[23][28] = 4'hA;
    SS1[24][28] = 4'hA;
    SS1[25][28] = 4'hD;
    SS1[26][28] = 4'hD;
    SS1[27][28] = 4'hC;
    SS1[28][28] = 4'hC;
    SS1[29][28] = 4'hD;
    SS1[30][28] = 4'hD;
    SS1[31][28] = 4'hD;
    SS1[32][28] = 4'hD;
    SS1[33][28] = 4'hD;
    SS1[34][28] = 4'hD;
    SS1[35][28] = 4'hD;
    SS1[36][28] = 4'hD;
    SS1[37][28] = 4'hD;
    SS1[38][28] = 4'h3;
    SS1[39][28] = 4'h3;
    SS1[40][28] = 4'h3;
    SS1[41][28] = 4'h0;
    SS1[42][28] = 4'h0;
    SS1[43][28] = 4'hD;
    SS1[44][28] = 4'hD;
    SS1[45][28] = 4'h0;
    SS1[46][28] = 4'h0;
    SS1[47][28] = 4'h0;
    SS1[0][29] = 4'h0;
    SS1[1][29] = 4'h0;
    SS1[2][29] = 4'h0;
    SS1[3][29] = 4'h0;
    SS1[4][29] = 4'h0;
    SS1[5][29] = 4'h0;
    SS1[6][29] = 4'h0;
    SS1[7][29] = 4'h0;
    SS1[8][29] = 4'h0;
    SS1[9][29] = 4'h0;
    SS1[10][29] = 4'h0;
    SS1[11][29] = 4'h0;
    SS1[12][29] = 4'h0;
    SS1[13][29] = 4'h0;
    SS1[14][29] = 4'h0;
    SS1[15][29] = 4'hC;
    SS1[16][29] = 4'hC;
    SS1[17][29] = 4'hC;
    SS1[18][29] = 4'hC;
    SS1[19][29] = 4'hC;
    SS1[20][29] = 4'hC;
    SS1[21][29] = 4'hC;
    SS1[22][29] = 4'hA;
    SS1[23][29] = 4'hA;
    SS1[24][29] = 4'hA;
    SS1[25][29] = 4'hD;
    SS1[26][29] = 4'hD;
    SS1[27][29] = 4'hD;
    SS1[28][29] = 4'hD;
    SS1[29][29] = 4'hD;
    SS1[30][29] = 4'hD;
    SS1[31][29] = 4'hD;
    SS1[32][29] = 4'hD;
    SS1[33][29] = 4'hD;
    SS1[34][29] = 4'hD;
    SS1[35][29] = 4'h0;
    SS1[36][29] = 4'h0;
    SS1[37][29] = 4'hD;
    SS1[38][29] = 4'h3;
    SS1[39][29] = 4'h3;
    SS1[40][29] = 4'h3;
    SS1[41][29] = 4'h0;
    SS1[42][29] = 4'h0;
    SS1[43][29] = 4'h0;
    SS1[44][29] = 4'h0;
    SS1[45][29] = 4'h0;
    SS1[46][29] = 4'h0;
    SS1[47][29] = 4'h0;
    SS1[0][30] = 4'h0;
    SS1[1][30] = 4'h0;
    SS1[2][30] = 4'h0;
    SS1[3][30] = 4'h0;
    SS1[4][30] = 4'h0;
    SS1[5][30] = 4'h0;
    SS1[6][30] = 4'h0;
    SS1[7][30] = 4'h0;
    SS1[8][30] = 4'h0;
    SS1[9][30] = 4'h0;
    SS1[10][30] = 4'h0;
    SS1[11][30] = 4'h0;
    SS1[12][30] = 4'h0;
    SS1[13][30] = 4'h0;
    SS1[14][30] = 4'h0;
    SS1[15][30] = 4'hD;
    SS1[16][30] = 4'hC;
    SS1[17][30] = 4'hC;
    SS1[18][30] = 4'hC;
    SS1[19][30] = 4'hC;
    SS1[20][30] = 4'hC;
    SS1[21][30] = 4'hC;
    SS1[22][30] = 4'hC;
    SS1[23][30] = 4'hC;
    SS1[24][30] = 4'hA;
    SS1[25][30] = 4'hD;
    SS1[26][30] = 4'hD;
    SS1[27][30] = 4'hD;
    SS1[28][30] = 4'hD;
    SS1[29][30] = 4'hD;
    SS1[30][30] = 4'hD;
    SS1[31][30] = 4'h3;
    SS1[32][30] = 4'hD;
    SS1[33][30] = 4'hD;
    SS1[34][30] = 4'h0;
    SS1[35][30] = 4'h0;
    SS1[36][30] = 4'h0;
    SS1[37][30] = 4'h0;
    SS1[38][30] = 4'h0;
    SS1[39][30] = 4'h0;
    SS1[40][30] = 4'h3;
    SS1[41][30] = 4'h0;
    SS1[42][30] = 4'h0;
    SS1[43][30] = 4'h0;
    SS1[44][30] = 4'h0;
    SS1[45][30] = 4'h0;
    SS1[46][30] = 4'h0;
    SS1[47][30] = 4'h0;
    SS1[0][31] = 4'h0;
    SS1[1][31] = 4'h0;
    SS1[2][31] = 4'h0;
    SS1[3][31] = 4'h0;
    SS1[4][31] = 4'h0;
    SS1[5][31] = 4'h0;
    SS1[6][31] = 4'h0;
    SS1[7][31] = 4'h0;
    SS1[8][31] = 4'h0;
    SS1[9][31] = 4'h0;
    SS1[10][31] = 4'h0;
    SS1[11][31] = 4'h0;
    SS1[12][31] = 4'h0;
    SS1[13][31] = 4'h0;
    SS1[14][31] = 4'hD;
    SS1[15][31] = 4'hD;
    SS1[16][31] = 4'hD;
    SS1[17][31] = 4'hD;
    SS1[18][31] = 4'hC;
    SS1[19][31] = 4'hC;
    SS1[20][31] = 4'hC;
    SS1[21][31] = 4'hC;
    SS1[22][31] = 4'hC;
    SS1[23][31] = 4'hC;
    SS1[24][31] = 4'hC;
    SS1[25][31] = 4'hC;
    SS1[26][31] = 4'hC;
    SS1[27][31] = 4'hD;
    SS1[28][31] = 4'hD;
    SS1[29][31] = 4'hD;
    SS1[30][31] = 4'hD;
    SS1[31][31] = 4'h3;
    SS1[32][31] = 4'h3;
    SS1[33][31] = 4'h3;
    SS1[34][31] = 4'h0;
    SS1[35][31] = 4'h0;
    SS1[36][31] = 4'h0;
    SS1[37][31] = 4'h0;
    SS1[38][31] = 4'h0;
    SS1[39][31] = 4'h0;
    SS1[40][31] = 4'h0;
    SS1[41][31] = 4'h0;
    SS1[42][31] = 4'h0;
    SS1[43][31] = 4'h0;
    SS1[44][31] = 4'h0;
    SS1[45][31] = 4'h0;
    SS1[46][31] = 4'h0;
    SS1[47][31] = 4'h0;
    SS1[0][32] = 4'h0;
    SS1[1][32] = 4'h0;
    SS1[2][32] = 4'h0;
    SS1[3][32] = 4'h0;
    SS1[4][32] = 4'h0;
    SS1[5][32] = 4'h0;
    SS1[6][32] = 4'h0;
    SS1[7][32] = 4'h0;
    SS1[8][32] = 4'h0;
    SS1[9][32] = 4'h0;
    SS1[10][32] = 4'h0;
    SS1[11][32] = 4'h0;
    SS1[12][32] = 4'h0;
    SS1[13][32] = 4'h0;
    SS1[14][32] = 4'hD;
    SS1[15][32] = 4'hD;
    SS1[16][32] = 4'hD;
    SS1[17][32] = 4'hC;
    SS1[18][32] = 4'hC;
    SS1[19][32] = 4'hC;
    SS1[20][32] = 4'hC;
    SS1[21][32] = 4'hC;
    SS1[22][32] = 4'hC;
    SS1[23][32] = 4'hC;
    SS1[24][32] = 4'hC;
    SS1[25][32] = 4'hC;
    SS1[26][32] = 4'hC;
    SS1[27][32] = 4'h0;
    SS1[28][32] = 4'h0;
    SS1[29][32] = 4'hD;
    SS1[30][32] = 4'h3;
    SS1[31][32] = 4'h3;
    SS1[32][32] = 4'h3;
    SS1[33][32] = 4'h0;
    SS1[34][32] = 4'h0;
    SS1[35][32] = 4'h0;
    SS1[36][32] = 4'h0;
    SS1[37][32] = 4'h0;
    SS1[38][32] = 4'h0;
    SS1[39][32] = 4'h0;
    SS1[40][32] = 4'h0;
    SS1[41][32] = 4'h0;
    SS1[42][32] = 4'h0;
    SS1[43][32] = 4'h0;
    SS1[44][32] = 4'h0;
    SS1[45][32] = 4'h0;
    SS1[46][32] = 4'h0;
    SS1[47][32] = 4'h0;
    SS1[0][33] = 4'h0;
    SS1[1][33] = 4'h0;
    SS1[2][33] = 4'h0;
    SS1[3][33] = 4'h0;
    SS1[4][33] = 4'h0;
    SS1[5][33] = 4'h0;
    SS1[6][33] = 4'h0;
    SS1[7][33] = 4'h0;
    SS1[8][33] = 4'h0;
    SS1[9][33] = 4'h0;
    SS1[10][33] = 4'h0;
    SS1[11][33] = 4'h0;
    SS1[12][33] = 4'h0;
    SS1[13][33] = 4'h0;
    SS1[14][33] = 4'hD;
    SS1[15][33] = 4'hD;
    SS1[16][33] = 4'hD;
    SS1[17][33] = 4'hC;
    SS1[18][33] = 4'hC;
    SS1[19][33] = 4'hC;
    SS1[20][33] = 4'hC;
    SS1[21][33] = 4'hC;
    SS1[22][33] = 4'hC;
    SS1[23][33] = 4'hD;
    SS1[24][33] = 4'hC;
    SS1[25][33] = 4'hC;
    SS1[26][33] = 4'hE;
    SS1[27][33] = 4'h0;
    SS1[28][33] = 4'h0;
    SS1[29][33] = 4'h0;
    SS1[30][33] = 4'h0;
    SS1[31][33] = 4'h3;
    SS1[32][33] = 4'h3;
    SS1[33][33] = 4'h0;
    SS1[34][33] = 4'h0;
    SS1[35][33] = 4'h0;
    SS1[36][33] = 4'h0;
    SS1[37][33] = 4'h0;
    SS1[38][33] = 4'h0;
    SS1[39][33] = 4'h0;
    SS1[40][33] = 4'h0;
    SS1[41][33] = 4'h0;
    SS1[42][33] = 4'h0;
    SS1[43][33] = 4'h0;
    SS1[44][33] = 4'h0;
    SS1[45][33] = 4'h0;
    SS1[46][33] = 4'h0;
    SS1[47][33] = 4'h0;
    SS1[0][34] = 4'h0;
    SS1[1][34] = 4'h0;
    SS1[2][34] = 4'h0;
    SS1[3][34] = 4'h0;
    SS1[4][34] = 4'h0;
    SS1[5][34] = 4'h0;
    SS1[6][34] = 4'h0;
    SS1[7][34] = 4'h0;
    SS1[8][34] = 4'h0;
    SS1[9][34] = 4'h0;
    SS1[10][34] = 4'h0;
    SS1[11][34] = 4'h0;
    SS1[12][34] = 4'h0;
    SS1[13][34] = 4'hD;
    SS1[14][34] = 4'hD;
    SS1[15][34] = 4'hD;
    SS1[16][34] = 4'hC;
    SS1[17][34] = 4'hC;
    SS1[18][34] = 4'hC;
    SS1[19][34] = 4'hC;
    SS1[20][34] = 4'hC;
    SS1[21][34] = 4'hC;
    SS1[22][34] = 4'hC;
    SS1[23][34] = 4'hD;
    SS1[24][34] = 4'hD;
    SS1[25][34] = 4'hD;
    SS1[26][34] = 4'h0;
    SS1[27][34] = 4'h0;
    SS1[28][34] = 4'h0;
    SS1[29][34] = 4'h0;
    SS1[30][34] = 4'h0;
    SS1[31][34] = 4'h0;
    SS1[32][34] = 4'h0;
    SS1[33][34] = 4'h0;
    SS1[34][34] = 4'h0;
    SS1[35][34] = 4'h0;
    SS1[36][34] = 4'h0;
    SS1[37][34] = 4'h0;
    SS1[38][34] = 4'h0;
    SS1[39][34] = 4'h0;
    SS1[40][34] = 4'h0;
    SS1[41][34] = 4'h0;
    SS1[42][34] = 4'h0;
    SS1[43][34] = 4'h0;
    SS1[44][34] = 4'h0;
    SS1[45][34] = 4'h0;
    SS1[46][34] = 4'h0;
    SS1[47][34] = 4'h0;
    SS1[0][35] = 4'h0;
    SS1[1][35] = 4'h0;
    SS1[2][35] = 4'h0;
    SS1[3][35] = 4'h0;
    SS1[4][35] = 4'h0;
    SS1[5][35] = 4'h0;
    SS1[6][35] = 4'h0;
    SS1[7][35] = 4'h0;
    SS1[8][35] = 4'h0;
    SS1[9][35] = 4'h0;
    SS1[10][35] = 4'h0;
    SS1[11][35] = 4'h0;
    SS1[12][35] = 4'h0;
    SS1[13][35] = 4'hD;
    SS1[14][35] = 4'hD;
    SS1[15][35] = 4'hD;
    SS1[16][35] = 4'hC;
    SS1[17][35] = 4'hC;
    SS1[18][35] = 4'hC;
    SS1[19][35] = 4'hC;
    SS1[20][35] = 4'hC;
    SS1[21][35] = 4'hC;
    SS1[22][35] = 4'hD;
    SS1[23][35] = 4'hD;
    SS1[24][35] = 4'hD;
    SS1[25][35] = 4'hD;
    SS1[26][35] = 4'h0;
    SS1[27][35] = 4'h0;
    SS1[28][35] = 4'h0;
    SS1[29][35] = 4'h0;
    SS1[30][35] = 4'h0;
    SS1[31][35] = 4'h0;
    SS1[32][35] = 4'h0;
    SS1[33][35] = 4'h0;
    SS1[34][35] = 4'h0;
    SS1[35][35] = 4'h0;
    SS1[36][35] = 4'h0;
    SS1[37][35] = 4'h0;
    SS1[38][35] = 4'h0;
    SS1[39][35] = 4'h0;
    SS1[40][35] = 4'h0;
    SS1[41][35] = 4'h0;
    SS1[42][35] = 4'h0;
    SS1[43][35] = 4'h0;
    SS1[44][35] = 4'h0;
    SS1[45][35] = 4'h0;
    SS1[46][35] = 4'h0;
    SS1[47][35] = 4'h0;
    SS1[0][36] = 4'h0;
    SS1[1][36] = 4'h0;
    SS1[2][36] = 4'h0;
    SS1[3][36] = 4'h0;
    SS1[4][36] = 4'h0;
    SS1[5][36] = 4'h0;
    SS1[6][36] = 4'h0;
    SS1[7][36] = 4'h0;
    SS1[8][36] = 4'h0;
    SS1[9][36] = 4'h0;
    SS1[10][36] = 4'h0;
    SS1[11][36] = 4'h0;
    SS1[12][36] = 4'hD;
    SS1[13][36] = 4'hD;
    SS1[14][36] = 4'hD;
    SS1[15][36] = 4'hD;
    SS1[16][36] = 4'hC;
    SS1[17][36] = 4'hC;
    SS1[18][36] = 4'hC;
    SS1[19][36] = 4'hC;
    SS1[20][36] = 4'hC;
    SS1[21][36] = 4'hC;
    SS1[22][36] = 4'hD;
    SS1[23][36] = 4'hD;
    SS1[24][36] = 4'hD;
    SS1[25][36] = 4'h0;
    SS1[26][36] = 4'h0;
    SS1[27][36] = 4'h0;
    SS1[28][36] = 4'h0;
    SS1[29][36] = 4'h0;
    SS1[30][36] = 4'h0;
    SS1[31][36] = 4'h0;
    SS1[32][36] = 4'h0;
    SS1[33][36] = 4'h0;
    SS1[34][36] = 4'h0;
    SS1[35][36] = 4'h0;
    SS1[36][36] = 4'h0;
    SS1[37][36] = 4'h0;
    SS1[38][36] = 4'h0;
    SS1[39][36] = 4'h0;
    SS1[40][36] = 4'h0;
    SS1[41][36] = 4'h0;
    SS1[42][36] = 4'h0;
    SS1[43][36] = 4'h0;
    SS1[44][36] = 4'h0;
    SS1[45][36] = 4'h0;
    SS1[46][36] = 4'h0;
    SS1[47][36] = 4'h0;
    SS1[0][37] = 4'h0;
    SS1[1][37] = 4'h0;
    SS1[2][37] = 4'h0;
    SS1[3][37] = 4'h0;
    SS1[4][37] = 4'h0;
    SS1[5][37] = 4'h0;
    SS1[6][37] = 4'h0;
    SS1[7][37] = 4'h0;
    SS1[8][37] = 4'h0;
    SS1[9][37] = 4'h0;
    SS1[10][37] = 4'h0;
    SS1[11][37] = 4'h0;
    SS1[12][37] = 4'hD;
    SS1[13][37] = 4'hD;
    SS1[14][37] = 4'hD;
    SS1[15][37] = 4'hC;
    SS1[16][37] = 4'hC;
    SS1[17][37] = 4'hC;
    SS1[18][37] = 4'hC;
    SS1[19][37] = 4'hC;
    SS1[20][37] = 4'hC;
    SS1[21][37] = 4'hC;
    SS1[22][37] = 4'hD;
    SS1[23][37] = 4'hD;
    SS1[24][37] = 4'hD;
    SS1[25][37] = 4'h0;
    SS1[26][37] = 4'h0;
    SS1[27][37] = 4'h0;
    SS1[28][37] = 4'h0;
    SS1[29][37] = 4'h0;
    SS1[30][37] = 4'h0;
    SS1[31][37] = 4'h0;
    SS1[32][37] = 4'h0;
    SS1[33][37] = 4'h0;
    SS1[34][37] = 4'h0;
    SS1[35][37] = 4'h0;
    SS1[36][37] = 4'h0;
    SS1[37][37] = 4'h0;
    SS1[38][37] = 4'h0;
    SS1[39][37] = 4'h0;
    SS1[40][37] = 4'h0;
    SS1[41][37] = 4'h0;
    SS1[42][37] = 4'h0;
    SS1[43][37] = 4'h0;
    SS1[44][37] = 4'h0;
    SS1[45][37] = 4'h0;
    SS1[46][37] = 4'h0;
    SS1[47][37] = 4'h0;
    SS1[0][38] = 4'h0;
    SS1[1][38] = 4'h0;
    SS1[2][38] = 4'h0;
    SS1[3][38] = 4'h0;
    SS1[4][38] = 4'h0;
    SS1[5][38] = 4'h0;
    SS1[6][38] = 4'h0;
    SS1[7][38] = 4'h0;
    SS1[8][38] = 4'h0;
    SS1[9][38] = 4'h0;
    SS1[10][38] = 4'h0;
    SS1[11][38] = 4'h0;
    SS1[12][38] = 4'hF;
    SS1[13][38] = 4'hD;
    SS1[14][38] = 4'hD;
    SS1[15][38] = 4'hC;
    SS1[16][38] = 4'hC;
    SS1[17][38] = 4'hC;
    SS1[18][38] = 4'hC;
    SS1[19][38] = 4'hC;
    SS1[20][38] = 4'hC;
    SS1[21][38] = 4'hD;
    SS1[22][38] = 4'hD;
    SS1[23][38] = 4'hD;
    SS1[24][38] = 4'h0;
    SS1[25][38] = 4'h0;
    SS1[26][38] = 4'h0;
    SS1[27][38] = 4'h0;
    SS1[28][38] = 4'h0;
    SS1[29][38] = 4'h0;
    SS1[30][38] = 4'h0;
    SS1[31][38] = 4'h0;
    SS1[32][38] = 4'h0;
    SS1[33][38] = 4'h0;
    SS1[34][38] = 4'h0;
    SS1[35][38] = 4'h0;
    SS1[36][38] = 4'h0;
    SS1[37][38] = 4'h0;
    SS1[38][38] = 4'h0;
    SS1[39][38] = 4'h0;
    SS1[40][38] = 4'h0;
    SS1[41][38] = 4'h0;
    SS1[42][38] = 4'h0;
    SS1[43][38] = 4'h0;
    SS1[44][38] = 4'h0;
    SS1[45][38] = 4'h0;
    SS1[46][38] = 4'h0;
    SS1[47][38] = 4'h0;
    SS1[0][39] = 4'h0;
    SS1[1][39] = 4'h0;
    SS1[2][39] = 4'h0;
    SS1[3][39] = 4'h0;
    SS1[4][39] = 4'h0;
    SS1[5][39] = 4'h0;
    SS1[6][39] = 4'h0;
    SS1[7][39] = 4'h0;
    SS1[8][39] = 4'h0;
    SS1[9][39] = 4'h0;
    SS1[10][39] = 4'h0;
    SS1[11][39] = 4'h0;
    SS1[12][39] = 4'h0;
    SS1[13][39] = 4'h0;
    SS1[14][39] = 4'hC;
    SS1[15][39] = 4'hC;
    SS1[16][39] = 4'hC;
    SS1[17][39] = 4'hC;
    SS1[18][39] = 4'hC;
    SS1[19][39] = 4'hC;
    SS1[20][39] = 4'hC;
    SS1[21][39] = 4'hD;
    SS1[22][39] = 4'hD;
    SS1[23][39] = 4'hD;
    SS1[24][39] = 4'h0;
    SS1[25][39] = 4'h0;
    SS1[26][39] = 4'h0;
    SS1[27][39] = 4'h0;
    SS1[28][39] = 4'h0;
    SS1[29][39] = 4'h0;
    SS1[30][39] = 4'h0;
    SS1[31][39] = 4'h0;
    SS1[32][39] = 4'h0;
    SS1[33][39] = 4'h0;
    SS1[34][39] = 4'h0;
    SS1[35][39] = 4'h0;
    SS1[36][39] = 4'h0;
    SS1[37][39] = 4'h0;
    SS1[38][39] = 4'h0;
    SS1[39][39] = 4'h0;
    SS1[40][39] = 4'h0;
    SS1[41][39] = 4'h0;
    SS1[42][39] = 4'h0;
    SS1[43][39] = 4'h0;
    SS1[44][39] = 4'h0;
    SS1[45][39] = 4'h0;
    SS1[46][39] = 4'h0;
    SS1[47][39] = 4'h0;
    SS1[0][40] = 4'h0;
    SS1[1][40] = 4'h0;
    SS1[2][40] = 4'h0;
    SS1[3][40] = 4'h0;
    SS1[4][40] = 4'h0;
    SS1[5][40] = 4'h0;
    SS1[6][40] = 4'h0;
    SS1[7][40] = 4'h0;
    SS1[8][40] = 4'h0;
    SS1[9][40] = 4'h0;
    SS1[10][40] = 4'h0;
    SS1[11][40] = 4'h0;
    SS1[12][40] = 4'h0;
    SS1[13][40] = 4'h0;
    SS1[14][40] = 4'hC;
    SS1[15][40] = 4'hC;
    SS1[16][40] = 4'hC;
    SS1[17][40] = 4'hC;
    SS1[18][40] = 4'hC;
    SS1[19][40] = 4'hC;
    SS1[20][40] = 4'hD;
    SS1[21][40] = 4'hD;
    SS1[22][40] = 4'hD;
    SS1[23][40] = 4'hD;
    SS1[24][40] = 4'h0;
    SS1[25][40] = 4'h0;
    SS1[26][40] = 4'h0;
    SS1[27][40] = 4'h0;
    SS1[28][40] = 4'h0;
    SS1[29][40] = 4'h0;
    SS1[30][40] = 4'h0;
    SS1[31][40] = 4'h0;
    SS1[32][40] = 4'h0;
    SS1[33][40] = 4'h0;
    SS1[34][40] = 4'h0;
    SS1[35][40] = 4'h0;
    SS1[36][40] = 4'h0;
    SS1[37][40] = 4'h0;
    SS1[38][40] = 4'h0;
    SS1[39][40] = 4'h0;
    SS1[40][40] = 4'h0;
    SS1[41][40] = 4'h0;
    SS1[42][40] = 4'h0;
    SS1[43][40] = 4'h0;
    SS1[44][40] = 4'h0;
    SS1[45][40] = 4'h0;
    SS1[46][40] = 4'h0;
    SS1[47][40] = 4'h0;
    SS1[0][41] = 4'h0;
    SS1[1][41] = 4'h0;
    SS1[2][41] = 4'h0;
    SS1[3][41] = 4'h0;
    SS1[4][41] = 4'h0;
    SS1[5][41] = 4'h0;
    SS1[6][41] = 4'h0;
    SS1[7][41] = 4'h0;
    SS1[8][41] = 4'h0;
    SS1[9][41] = 4'h0;
    SS1[10][41] = 4'h0;
    SS1[11][41] = 4'h0;
    SS1[12][41] = 4'h0;
    SS1[13][41] = 4'h0;
    SS1[14][41] = 4'hC;
    SS1[15][41] = 4'hC;
    SS1[16][41] = 4'hC;
    SS1[17][41] = 4'hC;
    SS1[18][41] = 4'hC;
    SS1[19][41] = 4'hC;
    SS1[20][41] = 4'hD;
    SS1[21][41] = 4'hD;
    SS1[22][41] = 4'hD;
    SS1[23][41] = 4'h0;
    SS1[24][41] = 4'h0;
    SS1[25][41] = 4'h0;
    SS1[26][41] = 4'h0;
    SS1[27][41] = 4'h0;
    SS1[28][41] = 4'h0;
    SS1[29][41] = 4'h0;
    SS1[30][41] = 4'h0;
    SS1[31][41] = 4'h0;
    SS1[32][41] = 4'h0;
    SS1[33][41] = 4'h0;
    SS1[34][41] = 4'h0;
    SS1[35][41] = 4'h0;
    SS1[36][41] = 4'h0;
    SS1[37][41] = 4'h0;
    SS1[38][41] = 4'h0;
    SS1[39][41] = 4'h0;
    SS1[40][41] = 4'h0;
    SS1[41][41] = 4'h0;
    SS1[42][41] = 4'h0;
    SS1[43][41] = 4'h0;
    SS1[44][41] = 4'h0;
    SS1[45][41] = 4'h0;
    SS1[46][41] = 4'h0;
    SS1[47][41] = 4'h0;
    SS1[0][42] = 4'h0;
    SS1[1][42] = 4'h0;
    SS1[2][42] = 4'h0;
    SS1[3][42] = 4'h0;
    SS1[4][42] = 4'h0;
    SS1[5][42] = 4'h0;
    SS1[6][42] = 4'h0;
    SS1[7][42] = 4'h0;
    SS1[8][42] = 4'h0;
    SS1[9][42] = 4'h0;
    SS1[10][42] = 4'h0;
    SS1[11][42] = 4'h0;
    SS1[12][42] = 4'h0;
    SS1[13][42] = 4'hC;
    SS1[14][42] = 4'hC;
    SS1[15][42] = 4'hC;
    SS1[16][42] = 4'hC;
    SS1[17][42] = 4'hC;
    SS1[18][42] = 4'hC;
    SS1[19][42] = 4'hC;
    SS1[20][42] = 4'h0;
    SS1[21][42] = 4'h0;
    SS1[22][42] = 4'hD;
    SS1[23][42] = 4'h0;
    SS1[24][42] = 4'h0;
    SS1[25][42] = 4'h0;
    SS1[26][42] = 4'h0;
    SS1[27][42] = 4'h0;
    SS1[28][42] = 4'h0;
    SS1[29][42] = 4'h0;
    SS1[30][42] = 4'h0;
    SS1[31][42] = 4'h0;
    SS1[32][42] = 4'h0;
    SS1[33][42] = 4'h0;
    SS1[34][42] = 4'h0;
    SS1[35][42] = 4'h0;
    SS1[36][42] = 4'h0;
    SS1[37][42] = 4'h0;
    SS1[38][42] = 4'h0;
    SS1[39][42] = 4'h0;
    SS1[40][42] = 4'h0;
    SS1[41][42] = 4'h0;
    SS1[42][42] = 4'h0;
    SS1[43][42] = 4'h0;
    SS1[44][42] = 4'h0;
    SS1[45][42] = 4'h0;
    SS1[46][42] = 4'h0;
    SS1[47][42] = 4'h0;
    SS1[0][43] = 4'h0;
    SS1[1][43] = 4'h0;
    SS1[2][43] = 4'h0;
    SS1[3][43] = 4'h0;
    SS1[4][43] = 4'h0;
    SS1[5][43] = 4'h0;
    SS1[6][43] = 4'h0;
    SS1[7][43] = 4'h0;
    SS1[8][43] = 4'h0;
    SS1[9][43] = 4'h0;
    SS1[10][43] = 4'h0;
    SS1[11][43] = 4'h0;
    SS1[12][43] = 4'h0;
    SS1[13][43] = 4'hC;
    SS1[14][43] = 4'hC;
    SS1[15][43] = 4'hC;
    SS1[16][43] = 4'hC;
    SS1[17][43] = 4'hC;
    SS1[18][43] = 4'hC;
    SS1[19][43] = 4'h0;
    SS1[20][43] = 4'h0;
    SS1[21][43] = 4'h0;
    SS1[22][43] = 4'h0;
    SS1[23][43] = 4'h0;
    SS1[24][43] = 4'h0;
    SS1[25][43] = 4'h0;
    SS1[26][43] = 4'h0;
    SS1[27][43] = 4'h0;
    SS1[28][43] = 4'h0;
    SS1[29][43] = 4'h0;
    SS1[30][43] = 4'h0;
    SS1[31][43] = 4'h0;
    SS1[32][43] = 4'h0;
    SS1[33][43] = 4'h0;
    SS1[34][43] = 4'h0;
    SS1[35][43] = 4'h0;
    SS1[36][43] = 4'h0;
    SS1[37][43] = 4'h0;
    SS1[38][43] = 4'h0;
    SS1[39][43] = 4'h0;
    SS1[40][43] = 4'h0;
    SS1[41][43] = 4'h0;
    SS1[42][43] = 4'h0;
    SS1[43][43] = 4'h0;
    SS1[44][43] = 4'h0;
    SS1[45][43] = 4'h0;
    SS1[46][43] = 4'h0;
    SS1[47][43] = 4'h0;
    SS1[0][44] = 4'h0;
    SS1[1][44] = 4'h0;
    SS1[2][44] = 4'h0;
    SS1[3][44] = 4'h0;
    SS1[4][44] = 4'h0;
    SS1[5][44] = 4'h0;
    SS1[6][44] = 4'h0;
    SS1[7][44] = 4'h0;
    SS1[8][44] = 4'h0;
    SS1[9][44] = 4'h0;
    SS1[10][44] = 4'h0;
    SS1[11][44] = 4'h0;
    SS1[12][44] = 4'hC;
    SS1[13][44] = 4'hC;
    SS1[14][44] = 4'hC;
    SS1[15][44] = 4'hC;
    SS1[16][44] = 4'hC;
    SS1[17][44] = 4'hC;
    SS1[18][44] = 4'hC;
    SS1[19][44] = 4'h0;
    SS1[20][44] = 4'h0;
    SS1[21][44] = 4'h0;
    SS1[22][44] = 4'h0;
    SS1[23][44] = 4'h0;
    SS1[24][44] = 4'h0;
    SS1[25][44] = 4'h0;
    SS1[26][44] = 4'h0;
    SS1[27][44] = 4'h0;
    SS1[28][44] = 4'h0;
    SS1[29][44] = 4'h0;
    SS1[30][44] = 4'h0;
    SS1[31][44] = 4'h0;
    SS1[32][44] = 4'h0;
    SS1[33][44] = 4'h0;
    SS1[34][44] = 4'h0;
    SS1[35][44] = 4'h0;
    SS1[36][44] = 4'h0;
    SS1[37][44] = 4'h0;
    SS1[38][44] = 4'h0;
    SS1[39][44] = 4'h0;
    SS1[40][44] = 4'h0;
    SS1[41][44] = 4'h0;
    SS1[42][44] = 4'h0;
    SS1[43][44] = 4'h0;
    SS1[44][44] = 4'h0;
    SS1[45][44] = 4'h0;
    SS1[46][44] = 4'h0;
    SS1[47][44] = 4'h0;
    SS1[0][45] = 4'h0;
    SS1[1][45] = 4'h0;
    SS1[2][45] = 4'h0;
    SS1[3][45] = 4'h0;
    SS1[4][45] = 4'h0;
    SS1[5][45] = 4'h0;
    SS1[6][45] = 4'h0;
    SS1[7][45] = 4'h0;
    SS1[8][45] = 4'h0;
    SS1[9][45] = 4'h0;
    SS1[10][45] = 4'h0;
    SS1[11][45] = 4'h0;
    SS1[12][45] = 4'h0;
    SS1[13][45] = 4'h0;
    SS1[14][45] = 4'hC;
    SS1[15][45] = 4'hC;
    SS1[16][45] = 4'hC;
    SS1[17][45] = 4'hC;
    SS1[18][45] = 4'h0;
    SS1[19][45] = 4'h0;
    SS1[20][45] = 4'h0;
    SS1[21][45] = 4'h0;
    SS1[22][45] = 4'h0;
    SS1[23][45] = 4'h0;
    SS1[24][45] = 4'h0;
    SS1[25][45] = 4'h0;
    SS1[26][45] = 4'h0;
    SS1[27][45] = 4'h0;
    SS1[28][45] = 4'h0;
    SS1[29][45] = 4'h0;
    SS1[30][45] = 4'h0;
    SS1[31][45] = 4'h0;
    SS1[32][45] = 4'h0;
    SS1[33][45] = 4'h0;
    SS1[34][45] = 4'h0;
    SS1[35][45] = 4'h0;
    SS1[36][45] = 4'h0;
    SS1[37][45] = 4'h0;
    SS1[38][45] = 4'h0;
    SS1[39][45] = 4'h0;
    SS1[40][45] = 4'h0;
    SS1[41][45] = 4'h0;
    SS1[42][45] = 4'h0;
    SS1[43][45] = 4'h0;
    SS1[44][45] = 4'h0;
    SS1[45][45] = 4'h0;
    SS1[46][45] = 4'h0;
    SS1[47][45] = 4'h0;
    SS1[0][46] = 4'h0;
    SS1[1][46] = 4'h0;
    SS1[2][46] = 4'h0;
    SS1[3][46] = 4'h0;
    SS1[4][46] = 4'h0;
    SS1[5][46] = 4'h0;
    SS1[6][46] = 4'h0;
    SS1[7][46] = 4'h0;
    SS1[8][46] = 4'h0;
    SS1[9][46] = 4'h0;
    SS1[10][46] = 4'h0;
    SS1[11][46] = 4'h0;
    SS1[12][46] = 4'h0;
    SS1[13][46] = 4'h0;
    SS1[14][46] = 4'h0;
    SS1[15][46] = 4'h0;
    SS1[16][46] = 4'hC;
    SS1[17][46] = 4'hC;
    SS1[18][46] = 4'h0;
    SS1[19][46] = 4'h0;
    SS1[20][46] = 4'h0;
    SS1[21][46] = 4'h0;
    SS1[22][46] = 4'h0;
    SS1[23][46] = 4'h0;
    SS1[24][46] = 4'h0;
    SS1[25][46] = 4'h0;
    SS1[26][46] = 4'h0;
    SS1[27][46] = 4'h0;
    SS1[28][46] = 4'h0;
    SS1[29][46] = 4'h0;
    SS1[30][46] = 4'h0;
    SS1[31][46] = 4'h0;
    SS1[32][46] = 4'h0;
    SS1[33][46] = 4'h0;
    SS1[34][46] = 4'h0;
    SS1[35][46] = 4'h0;
    SS1[36][46] = 4'h0;
    SS1[37][46] = 4'h0;
    SS1[38][46] = 4'h0;
    SS1[39][46] = 4'h0;
    SS1[40][46] = 4'h0;
    SS1[41][46] = 4'h0;
    SS1[42][46] = 4'h0;
    SS1[43][46] = 4'h0;
    SS1[44][46] = 4'h0;
    SS1[45][46] = 4'h0;
    SS1[46][46] = 4'h0;
    SS1[47][46] = 4'h0;
    SS1[0][47] = 4'h0;
    SS1[1][47] = 4'h0;
    SS1[2][47] = 4'h0;
    SS1[3][47] = 4'h0;
    SS1[4][47] = 4'h0;
    SS1[5][47] = 4'h0;
    SS1[6][47] = 4'h0;
    SS1[7][47] = 4'h0;
    SS1[8][47] = 4'h0;
    SS1[9][47] = 4'h0;
    SS1[10][47] = 4'h0;
    SS1[11][47] = 4'h0;
    SS1[12][47] = 4'h0;
    SS1[13][47] = 4'h0;
    SS1[14][47] = 4'h0;
    SS1[15][47] = 4'h0;
    SS1[16][47] = 4'h0;
    SS1[17][47] = 4'h0;
    SS1[18][47] = 4'h0;
    SS1[19][47] = 4'h0;
    SS1[20][47] = 4'h0;
    SS1[21][47] = 4'h0;
    SS1[22][47] = 4'h0;
    SS1[23][47] = 4'h0;
    SS1[24][47] = 4'h0;
    SS1[25][47] = 4'h0;
    SS1[26][47] = 4'h0;
    SS1[27][47] = 4'h0;
    SS1[28][47] = 4'h0;
    SS1[29][47] = 4'h0;
    SS1[30][47] = 4'h0;
    SS1[31][47] = 4'h0;
    SS1[32][47] = 4'h0;
    SS1[33][47] = 4'h0;
    SS1[34][47] = 4'h0;
    SS1[35][47] = 4'h0;
    SS1[36][47] = 4'h0;
    SS1[37][47] = 4'h0;
    SS1[38][47] = 4'h0;
    SS1[39][47] = 4'h0;
    SS1[40][47] = 4'h0;
    SS1[41][47] = 4'h0;
    SS1[42][47] = 4'h0;
    SS1[43][47] = 4'h0;
    SS1[44][47] = 4'h0;
    SS1[45][47] = 4'h0;
    SS1[46][47] = 4'h0;
    SS1[47][47] = 4'h0;
 
//SS 2
    SS2[0][0] = 4'h0;
    SS2[1][0] = 4'h0;
    SS2[2][0] = 4'h0;
    SS2[3][0] = 4'h0;
    SS2[4][0] = 4'h0;
    SS2[5][0] = 4'h0;
    SS2[6][0] = 4'h0;
    SS2[7][0] = 4'h0;
    SS2[8][0] = 4'h0;
    SS2[9][0] = 4'h0;
    SS2[10][0] = 4'h0;
    SS2[11][0] = 4'h0;
    SS2[12][0] = 4'h0;
    SS2[13][0] = 4'h0;
    SS2[14][0] = 4'h0;
    SS2[15][0] = 4'h0;
    SS2[16][0] = 4'h0;
    SS2[17][0] = 4'h0;
    SS2[18][0] = 4'h0;
    SS2[19][0] = 4'h0;
    SS2[20][0] = 4'h0;
    SS2[21][0] = 4'h0;
    SS2[22][0] = 4'h0;
    SS2[23][0] = 4'h0;
    SS2[24][0] = 4'h0;
    SS2[25][0] = 4'h0;
    SS2[26][0] = 4'h0;
    SS2[27][0] = 4'h0;
    SS2[28][0] = 4'h0;
    SS2[29][0] = 4'h0;
    SS2[30][0] = 4'h0;
    SS2[31][0] = 4'h0;
    SS2[32][0] = 4'h0;
    SS2[33][0] = 4'h0;
    SS2[34][0] = 4'h0;
    SS2[35][0] = 4'h0;
    SS2[36][0] = 4'h0;
    SS2[37][0] = 4'h0;
    SS2[38][0] = 4'h0;
    SS2[39][0] = 4'h0;
    SS2[40][0] = 4'h0;
    SS2[41][0] = 4'h0;
    SS2[42][0] = 4'h0;
    SS2[43][0] = 4'h0;
    SS2[44][0] = 4'h0;
    SS2[45][0] = 4'h0;
    SS2[46][0] = 4'h0;
    SS2[47][0] = 4'h0;
    SS2[0][1] = 4'h0;
    SS2[1][1] = 4'h0;
    SS2[2][1] = 4'h0;
    SS2[3][1] = 4'h0;
    SS2[4][1] = 4'h0;
    SS2[5][1] = 4'h0;
    SS2[6][1] = 4'h0;
    SS2[7][1] = 4'h0;
    SS2[8][1] = 4'h0;
    SS2[9][1] = 4'h0;
    SS2[10][1] = 4'h0;
    SS2[11][1] = 4'h0;
    SS2[12][1] = 4'h0;
    SS2[13][1] = 4'h0;
    SS2[14][1] = 4'h0;
    SS2[15][1] = 4'h0;
    SS2[16][1] = 4'h0;
    SS2[17][1] = 4'h0;
    SS2[18][1] = 4'h0;
    SS2[19][1] = 4'h0;
    SS2[20][1] = 4'h0;
    SS2[21][1] = 4'h0;
    SS2[22][1] = 4'h0;
    SS2[23][1] = 4'h0;
    SS2[24][1] = 4'h0;
    SS2[25][1] = 4'h0;
    SS2[26][1] = 4'h0;
    SS2[27][1] = 4'h0;
    SS2[28][1] = 4'h0;
    SS2[29][1] = 4'h0;
    SS2[30][1] = 4'h0;
    SS2[31][1] = 4'h0;
    SS2[32][1] = 4'h0;
    SS2[33][1] = 4'h0;
    SS2[34][1] = 4'h0;
    SS2[35][1] = 4'h0;
    SS2[36][1] = 4'h0;
    SS2[37][1] = 4'h0;
    SS2[38][1] = 4'h0;
    SS2[39][1] = 4'h0;
    SS2[40][1] = 4'h0;
    SS2[41][1] = 4'h0;
    SS2[42][1] = 4'h0;
    SS2[43][1] = 4'h0;
    SS2[44][1] = 4'h0;
    SS2[45][1] = 4'h0;
    SS2[46][1] = 4'h0;
    SS2[47][1] = 4'h0;
    SS2[0][2] = 4'h0;
    SS2[1][2] = 4'h0;
    SS2[2][2] = 4'h0;
    SS2[3][2] = 4'h0;
    SS2[4][2] = 4'h0;
    SS2[5][2] = 4'h0;
    SS2[6][2] = 4'h0;
    SS2[7][2] = 4'h0;
    SS2[8][2] = 4'h0;
    SS2[9][2] = 4'h0;
    SS2[10][2] = 4'h0;
    SS2[11][2] = 4'h0;
    SS2[12][2] = 4'h0;
    SS2[13][2] = 4'h0;
    SS2[14][2] = 4'h0;
    SS2[15][2] = 4'h0;
    SS2[16][2] = 4'h0;
    SS2[17][2] = 4'h0;
    SS2[18][2] = 4'h0;
    SS2[19][2] = 4'h0;
    SS2[20][2] = 4'h0;
    SS2[21][2] = 4'h0;
    SS2[22][2] = 4'h0;
    SS2[23][2] = 4'h0;
    SS2[24][2] = 4'h0;
    SS2[25][2] = 4'h0;
    SS2[26][2] = 4'h0;
    SS2[27][2] = 4'h0;
    SS2[28][2] = 4'h0;
    SS2[29][2] = 4'h0;
    SS2[30][2] = 4'h0;
    SS2[31][2] = 4'h0;
    SS2[32][2] = 4'h0;
    SS2[33][2] = 4'h0;
    SS2[34][2] = 4'h0;
    SS2[35][2] = 4'h0;
    SS2[36][2] = 4'h0;
    SS2[37][2] = 4'h0;
    SS2[38][2] = 4'h0;
    SS2[39][2] = 4'h0;
    SS2[40][2] = 4'h0;
    SS2[41][2] = 4'h0;
    SS2[42][2] = 4'h0;
    SS2[43][2] = 4'h0;
    SS2[44][2] = 4'h0;
    SS2[45][2] = 4'h0;
    SS2[46][2] = 4'h0;
    SS2[47][2] = 4'h0;
    SS2[0][3] = 4'h0;
    SS2[1][3] = 4'h0;
    SS2[2][3] = 4'h0;
    SS2[3][3] = 4'h0;
    SS2[4][3] = 4'h0;
    SS2[5][3] = 4'h0;
    SS2[6][3] = 4'h0;
    SS2[7][3] = 4'h0;
    SS2[8][3] = 4'h0;
    SS2[9][3] = 4'h0;
    SS2[10][3] = 4'h0;
    SS2[11][3] = 4'h0;
    SS2[12][3] = 4'h0;
    SS2[13][3] = 4'h0;
    SS2[14][3] = 4'h0;
    SS2[15][3] = 4'h0;
    SS2[16][3] = 4'h0;
    SS2[17][3] = 4'h0;
    SS2[18][3] = 4'h0;
    SS2[19][3] = 4'h0;
    SS2[20][3] = 4'h0;
    SS2[21][3] = 4'h0;
    SS2[22][3] = 4'h0;
    SS2[23][3] = 4'h0;
    SS2[24][3] = 4'h0;
    SS2[25][3] = 4'h0;
    SS2[26][3] = 4'h0;
    SS2[27][3] = 4'h0;
    SS2[28][3] = 4'h0;
    SS2[29][3] = 4'h0;
    SS2[30][3] = 4'h0;
    SS2[31][3] = 4'h0;
    SS2[32][3] = 4'h0;
    SS2[33][3] = 4'h0;
    SS2[34][3] = 4'h0;
    SS2[35][3] = 4'h0;
    SS2[36][3] = 4'h0;
    SS2[37][3] = 4'h0;
    SS2[38][3] = 4'h0;
    SS2[39][3] = 4'h0;
    SS2[40][3] = 4'h0;
    SS2[41][3] = 4'h0;
    SS2[42][3] = 4'h0;
    SS2[43][3] = 4'h0;
    SS2[44][3] = 4'h0;
    SS2[45][3] = 4'h0;
    SS2[46][3] = 4'h0;
    SS2[47][3] = 4'h0;
    SS2[0][4] = 4'h0;
    SS2[1][4] = 4'h0;
    SS2[2][4] = 4'h0;
    SS2[3][4] = 4'h0;
    SS2[4][4] = 4'h0;
    SS2[5][4] = 4'h0;
    SS2[6][4] = 4'h0;
    SS2[7][4] = 4'h0;
    SS2[8][4] = 4'h0;
    SS2[9][4] = 4'h0;
    SS2[10][4] = 4'h0;
    SS2[11][4] = 4'h0;
    SS2[12][4] = 4'h0;
    SS2[13][4] = 4'h0;
    SS2[14][4] = 4'h0;
    SS2[15][4] = 4'h0;
    SS2[16][4] = 4'h0;
    SS2[17][4] = 4'h0;
    SS2[18][4] = 4'h0;
    SS2[19][4] = 4'h0;
    SS2[20][4] = 4'h0;
    SS2[21][4] = 4'h0;
    SS2[22][4] = 4'h0;
    SS2[23][4] = 4'h0;
    SS2[24][4] = 4'h0;
    SS2[25][4] = 4'h0;
    SS2[26][4] = 4'h0;
    SS2[27][4] = 4'h0;
    SS2[28][4] = 4'h0;
    SS2[29][4] = 4'h0;
    SS2[30][4] = 4'h0;
    SS2[31][4] = 4'h0;
    SS2[32][4] = 4'h0;
    SS2[33][4] = 4'h0;
    SS2[34][4] = 4'h0;
    SS2[35][4] = 4'h0;
    SS2[36][4] = 4'h0;
    SS2[37][4] = 4'h0;
    SS2[38][4] = 4'h0;
    SS2[39][4] = 4'h0;
    SS2[40][4] = 4'h0;
    SS2[41][4] = 4'h0;
    SS2[42][4] = 4'h0;
    SS2[43][4] = 4'h0;
    SS2[44][4] = 4'h0;
    SS2[45][4] = 4'h0;
    SS2[46][4] = 4'h0;
    SS2[47][4] = 4'h0;
    SS2[0][5] = 4'h0;
    SS2[1][5] = 4'h0;
    SS2[2][5] = 4'h0;
    SS2[3][5] = 4'h0;
    SS2[4][5] = 4'h0;
    SS2[5][5] = 4'h0;
    SS2[6][5] = 4'h0;
    SS2[7][5] = 4'h0;
    SS2[8][5] = 4'h0;
    SS2[9][5] = 4'h0;
    SS2[10][5] = 4'h0;
    SS2[11][5] = 4'h0;
    SS2[12][5] = 4'h0;
    SS2[13][5] = 4'h0;
    SS2[14][5] = 4'h0;
    SS2[15][5] = 4'h0;
    SS2[16][5] = 4'h0;
    SS2[17][5] = 4'h0;
    SS2[18][5] = 4'h0;
    SS2[19][5] = 4'h0;
    SS2[20][5] = 4'h0;
    SS2[21][5] = 4'h0;
    SS2[22][5] = 4'h0;
    SS2[23][5] = 4'h0;
    SS2[24][5] = 4'h0;
    SS2[25][5] = 4'h0;
    SS2[26][5] = 4'h0;
    SS2[27][5] = 4'h0;
    SS2[28][5] = 4'h0;
    SS2[29][5] = 4'h0;
    SS2[30][5] = 4'h0;
    SS2[31][5] = 4'h0;
    SS2[32][5] = 4'h0;
    SS2[33][5] = 4'h0;
    SS2[34][5] = 4'h0;
    SS2[35][5] = 4'h0;
    SS2[36][5] = 4'h0;
    SS2[37][5] = 4'h0;
    SS2[38][5] = 4'hC;
    SS2[39][5] = 4'h0;
    SS2[40][5] = 4'h0;
    SS2[41][5] = 4'h0;
    SS2[42][5] = 4'h0;
    SS2[43][5] = 4'h0;
    SS2[44][5] = 4'h0;
    SS2[45][5] = 4'h0;
    SS2[46][5] = 4'h0;
    SS2[47][5] = 4'h0;
    SS2[0][6] = 4'h0;
    SS2[1][6] = 4'h0;
    SS2[2][6] = 4'h0;
    SS2[3][6] = 4'h0;
    SS2[4][6] = 4'h0;
    SS2[5][6] = 4'h0;
    SS2[6][6] = 4'h0;
    SS2[7][6] = 4'h0;
    SS2[8][6] = 4'h0;
    SS2[9][6] = 4'h0;
    SS2[10][6] = 4'h0;
    SS2[11][6] = 4'h0;
    SS2[12][6] = 4'h0;
    SS2[13][6] = 4'h0;
    SS2[14][6] = 4'h0;
    SS2[15][6] = 4'h0;
    SS2[16][6] = 4'h0;
    SS2[17][6] = 4'h0;
    SS2[18][6] = 4'h0;
    SS2[19][6] = 4'h0;
    SS2[20][6] = 4'h0;
    SS2[21][6] = 4'h0;
    SS2[22][6] = 4'h0;
    SS2[23][6] = 4'h0;
    SS2[24][6] = 4'h0;
    SS2[25][6] = 4'h0;
    SS2[26][6] = 4'h0;
    SS2[27][6] = 4'h0;
    SS2[28][6] = 4'h0;
    SS2[29][6] = 4'h0;
    SS2[30][6] = 4'h0;
    SS2[31][6] = 4'h0;
    SS2[32][6] = 4'h0;
    SS2[33][6] = 4'h0;
    SS2[34][6] = 4'h0;
    SS2[35][6] = 4'h0;
    SS2[36][6] = 4'h0;
    SS2[37][6] = 4'hC;
    SS2[38][6] = 4'hC;
    SS2[39][6] = 4'hC;
    SS2[40][6] = 4'h0;
    SS2[41][6] = 4'h0;
    SS2[42][6] = 4'h0;
    SS2[43][6] = 4'h0;
    SS2[44][6] = 4'h0;
    SS2[45][6] = 4'h0;
    SS2[46][6] = 4'h0;
    SS2[47][6] = 4'h0;
    SS2[0][7] = 4'h0;
    SS2[1][7] = 4'h0;
    SS2[2][7] = 4'h0;
    SS2[3][7] = 4'h0;
    SS2[4][7] = 4'h0;
    SS2[5][7] = 4'h0;
    SS2[6][7] = 4'h0;
    SS2[7][7] = 4'h0;
    SS2[8][7] = 4'h0;
    SS2[9][7] = 4'h0;
    SS2[10][7] = 4'h0;
    SS2[11][7] = 4'h0;
    SS2[12][7] = 4'h0;
    SS2[13][7] = 4'h0;
    SS2[14][7] = 4'h0;
    SS2[15][7] = 4'h0;
    SS2[16][7] = 4'h0;
    SS2[17][7] = 4'h0;
    SS2[18][7] = 4'h0;
    SS2[19][7] = 4'h0;
    SS2[20][7] = 4'h0;
    SS2[21][7] = 4'h0;
    SS2[22][7] = 4'h0;
    SS2[23][7] = 4'h0;
    SS2[24][7] = 4'h0;
    SS2[25][7] = 4'h0;
    SS2[26][7] = 4'h0;
    SS2[27][7] = 4'h0;
    SS2[28][7] = 4'h0;
    SS2[29][7] = 4'h0;
    SS2[30][7] = 4'h0;
    SS2[31][7] = 4'h0;
    SS2[32][7] = 4'hD;
    SS2[33][7] = 4'h0;
    SS2[34][7] = 4'h0;
    SS2[35][7] = 4'h0;
    SS2[36][7] = 4'hC;
    SS2[37][7] = 4'hC;
    SS2[38][7] = 4'hC;
    SS2[39][7] = 4'hC;
    SS2[40][7] = 4'hC;
    SS2[41][7] = 4'h0;
    SS2[42][7] = 4'h0;
    SS2[43][7] = 4'h0;
    SS2[44][7] = 4'h0;
    SS2[45][7] = 4'h0;
    SS2[46][7] = 4'h0;
    SS2[47][7] = 4'h0;
    SS2[0][8] = 4'h0;
    SS2[1][8] = 4'h0;
    SS2[2][8] = 4'h0;
    SS2[3][8] = 4'h0;
    SS2[4][8] = 4'h0;
    SS2[5][8] = 4'h0;
    SS2[6][8] = 4'h0;
    SS2[7][8] = 4'h0;
    SS2[8][8] = 4'h0;
    SS2[9][8] = 4'h0;
    SS2[10][8] = 4'h0;
    SS2[11][8] = 4'h0;
    SS2[12][8] = 4'h0;
    SS2[13][8] = 4'h0;
    SS2[14][8] = 4'h0;
    SS2[15][8] = 4'h0;
    SS2[16][8] = 4'h0;
    SS2[17][8] = 4'h0;
    SS2[18][8] = 4'h0;
    SS2[19][8] = 4'h0;
    SS2[20][8] = 4'h0;
    SS2[21][8] = 4'h0;
    SS2[22][8] = 4'h0;
    SS2[23][8] = 4'h0;
    SS2[24][8] = 4'h0;
    SS2[25][8] = 4'h0;
    SS2[26][8] = 4'h0;
    SS2[27][8] = 4'h0;
    SS2[28][8] = 4'h0;
    SS2[29][8] = 4'h0;
    SS2[30][8] = 4'h0;
    SS2[31][8] = 4'hD;
    SS2[32][8] = 4'hD;
    SS2[33][8] = 4'hD;
    SS2[34][8] = 4'h0;
    SS2[35][8] = 4'hC;
    SS2[36][8] = 4'hC;
    SS2[37][8] = 4'hC;
    SS2[38][8] = 4'hC;
    SS2[39][8] = 4'hC;
    SS2[40][8] = 4'hC;
    SS2[41][8] = 4'hC;
    SS2[42][8] = 4'h0;
    SS2[43][8] = 4'h0;
    SS2[44][8] = 4'h0;
    SS2[45][8] = 4'h0;
    SS2[46][8] = 4'h0;
    SS2[47][8] = 4'h0;
    SS2[0][9] = 4'h0;
    SS2[1][9] = 4'h0;
    SS2[2][9] = 4'h0;
    SS2[3][9] = 4'h0;
    SS2[4][9] = 4'h0;
    SS2[5][9] = 4'h0;
    SS2[6][9] = 4'h0;
    SS2[7][9] = 4'h0;
    SS2[8][9] = 4'h0;
    SS2[9][9] = 4'h0;
    SS2[10][9] = 4'h0;
    SS2[11][9] = 4'h0;
    SS2[12][9] = 4'h0;
    SS2[13][9] = 4'h0;
    SS2[14][9] = 4'h0;
    SS2[15][9] = 4'h0;
    SS2[16][9] = 4'h0;
    SS2[17][9] = 4'h0;
    SS2[18][9] = 4'h0;
    SS2[19][9] = 4'h0;
    SS2[20][9] = 4'h0;
    SS2[21][9] = 4'h0;
    SS2[22][9] = 4'h0;
    SS2[23][9] = 4'h0;
    SS2[24][9] = 4'h0;
    SS2[25][9] = 4'h0;
    SS2[26][9] = 4'h0;
    SS2[27][9] = 4'h0;
    SS2[28][9] = 4'h0;
    SS2[29][9] = 4'h0;
    SS2[30][9] = 4'hD;
    SS2[31][9] = 4'hD;
    SS2[32][9] = 4'hD;
    SS2[33][9] = 4'hD;
    SS2[34][9] = 4'hC;
    SS2[35][9] = 4'hC;
    SS2[36][9] = 4'hC;
    SS2[37][9] = 4'hC;
    SS2[38][9] = 4'hC;
    SS2[39][9] = 4'hC;
    SS2[40][9] = 4'hC;
    SS2[41][9] = 4'hC;
    SS2[42][9] = 4'hC;
    SS2[43][9] = 4'h0;
    SS2[44][9] = 4'h0;
    SS2[45][9] = 4'h0;
    SS2[46][9] = 4'h0;
    SS2[47][9] = 4'h0;
    SS2[0][10] = 4'h0;
    SS2[1][10] = 4'h0;
    SS2[2][10] = 4'h0;
    SS2[3][10] = 4'h0;
    SS2[4][10] = 4'h0;
    SS2[5][10] = 4'h0;
    SS2[6][10] = 4'h0;
    SS2[7][10] = 4'h0;
    SS2[8][10] = 4'h0;
    SS2[9][10] = 4'h0;
    SS2[10][10] = 4'h0;
    SS2[11][10] = 4'h0;
    SS2[12][10] = 4'h0;
    SS2[13][10] = 4'h0;
    SS2[14][10] = 4'h0;
    SS2[15][10] = 4'h0;
    SS2[16][10] = 4'h0;
    SS2[17][10] = 4'h0;
    SS2[18][10] = 4'h0;
    SS2[19][10] = 4'h0;
    SS2[20][10] = 4'h0;
    SS2[21][10] = 4'h0;
    SS2[22][10] = 4'h0;
    SS2[23][10] = 4'h0;
    SS2[24][10] = 4'h0;
    SS2[25][10] = 4'h0;
    SS2[26][10] = 4'h0;
    SS2[27][10] = 4'h0;
    SS2[28][10] = 4'h0;
    SS2[29][10] = 4'hD;
    SS2[30][10] = 4'hD;
    SS2[31][10] = 4'hD;
    SS2[32][10] = 4'hD;
    SS2[33][10] = 4'hC;
    SS2[34][10] = 4'hC;
    SS2[35][10] = 4'hC;
    SS2[36][10] = 4'hC;
    SS2[37][10] = 4'hC;
    SS2[38][10] = 4'hC;
    SS2[39][10] = 4'hC;
    SS2[40][10] = 4'hC;
    SS2[41][10] = 4'hC;
    SS2[42][10] = 4'h0;
    SS2[43][10] = 4'h0;
    SS2[44][10] = 4'h0;
    SS2[45][10] = 4'h0;
    SS2[46][10] = 4'h0;
    SS2[47][10] = 4'h0;
    SS2[0][11] = 4'h0;
    SS2[1][11] = 4'h0;
    SS2[2][11] = 4'h0;
    SS2[3][11] = 4'h0;
    SS2[4][11] = 4'h0;
    SS2[5][11] = 4'h0;
    SS2[6][11] = 4'h0;
    SS2[7][11] = 4'h0;
    SS2[8][11] = 4'h0;
    SS2[9][11] = 4'h0;
    SS2[10][11] = 4'h0;
    SS2[11][11] = 4'h2;
    SS2[12][11] = 4'h0;
    SS2[13][11] = 4'h0;
    SS2[14][11] = 4'h0;
    SS2[15][11] = 4'h0;
    SS2[16][11] = 4'h0;
    SS2[17][11] = 4'h0;
    SS2[18][11] = 4'h0;
    SS2[19][11] = 4'h2;
    SS2[20][11] = 4'h0;
    SS2[21][11] = 4'h0;
    SS2[22][11] = 4'h0;
    SS2[23][11] = 4'h0;
    SS2[24][11] = 4'h0;
    SS2[25][11] = 4'h0;
    SS2[26][11] = 4'h0;
    SS2[27][11] = 4'h0;
    SS2[28][11] = 4'hD;
    SS2[29][11] = 4'hD;
    SS2[30][11] = 4'hD;
    SS2[31][11] = 4'hD;
    SS2[32][11] = 4'hC;
    SS2[33][11] = 4'hC;
    SS2[34][11] = 4'hC;
    SS2[35][11] = 4'hC;
    SS2[36][11] = 4'hC;
    SS2[37][11] = 4'hC;
    SS2[38][11] = 4'hC;
    SS2[39][11] = 4'hC;
    SS2[40][11] = 4'hC;
    SS2[41][11] = 4'h0;
    SS2[42][11] = 4'h0;
    SS2[43][11] = 4'h0;
    SS2[44][11] = 4'h0;
    SS2[45][11] = 4'h0;
    SS2[46][11] = 4'h0;
    SS2[47][11] = 4'h0;
    SS2[0][12] = 4'h0;
    SS2[1][12] = 4'h0;
    SS2[2][12] = 4'hD;
    SS2[3][12] = 4'hD;
    SS2[4][12] = 4'h0;
    SS2[5][12] = 4'h0;
    SS2[6][12] = 4'hD;
    SS2[7][12] = 4'hD;
    SS2[8][12] = 4'h0;
    SS2[9][12] = 4'h0;
    SS2[10][12] = 4'h3;
    SS2[11][12] = 4'h3;
    SS2[12][12] = 4'h2;
    SS2[13][12] = 4'h0;
    SS2[14][12] = 4'h0;
    SS2[15][12] = 4'h0;
    SS2[16][12] = 4'h0;
    SS2[17][12] = 4'h0;
    SS2[18][12] = 4'h2;
    SS2[19][12] = 4'h3;
    SS2[20][12] = 4'h3;
    SS2[21][12] = 4'h0;
    SS2[22][12] = 4'h0;
    SS2[23][12] = 4'h0;
    SS2[24][12] = 4'h0;
    SS2[25][12] = 4'h0;
    SS2[26][12] = 4'h0;
    SS2[27][12] = 4'hD;
    SS2[28][12] = 4'hD;
    SS2[29][12] = 4'hD;
    SS2[30][12] = 4'hD;
    SS2[31][12] = 4'hC;
    SS2[32][12] = 4'hC;
    SS2[33][12] = 4'hC;
    SS2[34][12] = 4'hC;
    SS2[35][12] = 4'hC;
    SS2[36][12] = 4'hC;
    SS2[37][12] = 4'hC;
    SS2[38][12] = 4'hC;
    SS2[39][12] = 4'hC;
    SS2[40][12] = 4'h0;
    SS2[41][12] = 4'h0;
    SS2[42][12] = 4'h0;
    SS2[43][12] = 4'h0;
    SS2[44][12] = 4'h0;
    SS2[45][12] = 4'h0;
    SS2[46][12] = 4'h0;
    SS2[47][12] = 4'h0;
    SS2[0][13] = 4'h0;
    SS2[1][13] = 4'hD;
    SS2[2][13] = 4'hD;
    SS2[3][13] = 4'hD;
    SS2[4][13] = 4'hD;
    SS2[5][13] = 4'hD;
    SS2[6][13] = 4'hD;
    SS2[7][13] = 4'hD;
    SS2[8][13] = 4'hD;
    SS2[9][13] = 4'h3;
    SS2[10][13] = 4'h3;
    SS2[11][13] = 4'h3;
    SS2[12][13] = 4'h3;
    SS2[13][13] = 4'hE;
    SS2[14][13] = 4'h0;
    SS2[15][13] = 4'h0;
    SS2[16][13] = 4'h0;
    SS2[17][13] = 4'h0;
    SS2[18][13] = 4'h3;
    SS2[19][13] = 4'h3;
    SS2[20][13] = 4'h3;
    SS2[21][13] = 4'h3;
    SS2[22][13] = 4'h0;
    SS2[23][13] = 4'h0;
    SS2[24][13] = 4'h0;
    SS2[25][13] = 4'h0;
    SS2[26][13] = 4'hD;
    SS2[27][13] = 4'hD;
    SS2[28][13] = 4'hD;
    SS2[29][13] = 4'hD;
    SS2[30][13] = 4'hC;
    SS2[31][13] = 4'hC;
    SS2[32][13] = 4'hC;
    SS2[33][13] = 4'hC;
    SS2[34][13] = 4'hC;
    SS2[35][13] = 4'hC;
    SS2[36][13] = 4'hC;
    SS2[37][13] = 4'hC;
    SS2[38][13] = 4'hC;
    SS2[39][13] = 4'h0;
    SS2[40][13] = 4'h0;
    SS2[41][13] = 4'h0;
    SS2[42][13] = 4'h0;
    SS2[43][13] = 4'h0;
    SS2[44][13] = 4'h0;
    SS2[45][13] = 4'h0;
    SS2[46][13] = 4'h0;
    SS2[47][13] = 4'h0;
    SS2[0][14] = 4'h0;
    SS2[1][14] = 4'h0;
    SS2[2][14] = 4'hD;
    SS2[3][14] = 4'hD;
    SS2[4][14] = 4'hD;
    SS2[5][14] = 4'hD;
    SS2[6][14] = 4'hD;
    SS2[7][14] = 4'hD;
    SS2[8][14] = 4'hD;
    SS2[9][14] = 4'hD;
    SS2[10][14] = 4'h3;
    SS2[11][14] = 4'h3;
    SS2[12][14] = 4'hD;
    SS2[13][14] = 4'hD;
    SS2[14][14] = 4'hE;
    SS2[15][14] = 4'h0;
    SS2[16][14] = 4'h0;
    SS2[17][14] = 4'hD;
    SS2[18][14] = 4'hD;
    SS2[19][14] = 4'h3;
    SS2[20][14] = 4'h3;
    SS2[21][14] = 4'hD;
    SS2[22][14] = 4'hD;
    SS2[23][14] = 4'h0;
    SS2[24][14] = 4'h0;
    SS2[25][14] = 4'hC;
    SS2[26][14] = 4'hC;
    SS2[27][14] = 4'hD;
    SS2[28][14] = 4'hD;
    SS2[29][14] = 4'hC;
    SS2[30][14] = 4'hC;
    SS2[31][14] = 4'hC;
    SS2[32][14] = 4'hC;
    SS2[33][14] = 4'hC;
    SS2[34][14] = 4'hC;
    SS2[35][14] = 4'hC;
    SS2[36][14] = 4'hC;
    SS2[37][14] = 4'hC;
    SS2[38][14] = 4'hD;
    SS2[39][14] = 4'hD;
    SS2[40][14] = 4'h0;
    SS2[41][14] = 4'h0;
    SS2[42][14] = 4'h0;
    SS2[43][14] = 4'h0;
    SS2[44][14] = 4'h0;
    SS2[45][14] = 4'h0;
    SS2[46][14] = 4'h0;
    SS2[47][14] = 4'h0;
    SS2[0][15] = 4'h0;
    SS2[1][15] = 4'h0;
    SS2[2][15] = 4'h0;
    SS2[3][15] = 4'hD;
    SS2[4][15] = 4'hD;
    SS2[5][15] = 4'hD;
    SS2[6][15] = 4'hD;
    SS2[7][15] = 4'hD;
    SS2[8][15] = 4'hD;
    SS2[9][15] = 4'hD;
    SS2[10][15] = 4'hD;
    SS2[11][15] = 4'hD;
    SS2[12][15] = 4'hD;
    SS2[13][15] = 4'hD;
    SS2[14][15] = 4'hD;
    SS2[15][15] = 4'hD;
    SS2[16][15] = 4'hD;
    SS2[17][15] = 4'hD;
    SS2[18][15] = 4'hD;
    SS2[19][15] = 4'hD;
    SS2[20][15] = 4'hD;
    SS2[21][15] = 4'hD;
    SS2[22][15] = 4'hD;
    SS2[23][15] = 4'hD;
    SS2[24][15] = 4'hC;
    SS2[25][15] = 4'hC;
    SS2[26][15] = 4'hC;
    SS2[27][15] = 4'hC;
    SS2[28][15] = 4'hC;
    SS2[29][15] = 4'hC;
    SS2[30][15] = 4'hC;
    SS2[31][15] = 4'hC;
    SS2[32][15] = 4'hC;
    SS2[33][15] = 4'hC;
    SS2[34][15] = 4'hC;
    SS2[35][15] = 4'hC;
    SS2[36][15] = 4'hC;
    SS2[37][15] = 4'hD;
    SS2[38][15] = 4'hD;
    SS2[39][15] = 4'hD;
    SS2[40][15] = 4'hD;
    SS2[41][15] = 4'h0;
    SS2[42][15] = 4'h0;
    SS2[43][15] = 4'h0;
    SS2[44][15] = 4'h0;
    SS2[45][15] = 4'h0;
    SS2[46][15] = 4'h0;
    SS2[47][15] = 4'h0;
    SS2[0][16] = 4'h0;
    SS2[1][16] = 4'h0;
    SS2[2][16] = 4'h0;
    SS2[3][16] = 4'h0;
    SS2[4][16] = 4'hD;
    SS2[5][16] = 4'hD;
    SS2[6][16] = 4'hE;
    SS2[7][16] = 4'hE;
    SS2[8][16] = 4'hD;
    SS2[9][16] = 4'hD;
    SS2[10][16] = 4'hE;
    SS2[11][16] = 4'hE;
    SS2[12][16] = 4'hD;
    SS2[13][16] = 4'hD;
    SS2[14][16] = 4'hD;
    SS2[15][16] = 4'hD;
    SS2[16][16] = 4'hD;
    SS2[17][16] = 4'hD;
    SS2[18][16] = 4'hD;
    SS2[19][16] = 4'hD;
    SS2[20][16] = 4'hD;
    SS2[21][16] = 4'hD;
    SS2[22][16] = 4'hD;
    SS2[23][16] = 4'hD;
    SS2[24][16] = 4'hD;
    SS2[25][16] = 4'hC;
    SS2[26][16] = 4'hC;
    SS2[27][16] = 4'hC;
    SS2[28][16] = 4'hC;
    SS2[29][16] = 4'hC;
    SS2[30][16] = 4'hC;
    SS2[31][16] = 4'hC;
    SS2[32][16] = 4'hC;
    SS2[33][16] = 4'hC;
    SS2[34][16] = 4'hC;
    SS2[35][16] = 4'hC;
    SS2[36][16] = 4'hD;
    SS2[37][16] = 4'hD;
    SS2[38][16] = 4'hD;
    SS2[39][16] = 4'hD;
    SS2[40][16] = 4'h0;
    SS2[41][16] = 4'h0;
    SS2[42][16] = 4'h0;
    SS2[43][16] = 4'h0;
    SS2[44][16] = 4'h0;
    SS2[45][16] = 4'h0;
    SS2[46][16] = 4'h0;
    SS2[47][16] = 4'h0;
    SS2[0][17] = 4'h0;
    SS2[1][17] = 4'h0;
    SS2[2][17] = 4'h0;
    SS2[3][17] = 4'h0;
    SS2[4][17] = 4'h0;
    SS2[5][17] = 4'hE;
    SS2[6][17] = 4'hE;
    SS2[7][17] = 4'hE;
    SS2[8][17] = 4'hE;
    SS2[9][17] = 4'hE;
    SS2[10][17] = 4'hE;
    SS2[11][17] = 4'hE;
    SS2[12][17] = 4'hE;
    SS2[13][17] = 4'hD;
    SS2[14][17] = 4'hD;
    SS2[15][17] = 4'hD;
    SS2[16][17] = 4'hD;
    SS2[17][17] = 4'hD;
    SS2[18][17] = 4'hD;
    SS2[19][17] = 4'hD;
    SS2[20][17] = 4'hD;
    SS2[21][17] = 4'hD;
    SS2[22][17] = 4'hD;
    SS2[23][17] = 4'hD;
    SS2[24][17] = 4'hD;
    SS2[25][17] = 4'hD;
    SS2[26][17] = 4'hC;
    SS2[27][17] = 4'hC;
    SS2[28][17] = 4'hC;
    SS2[29][17] = 4'hC;
    SS2[30][17] = 4'hC;
    SS2[31][17] = 4'hC;
    SS2[32][17] = 4'hC;
    SS2[33][17] = 4'hC;
    SS2[34][17] = 4'hC;
    SS2[35][17] = 4'hD;
    SS2[36][17] = 4'hD;
    SS2[37][17] = 4'hD;
    SS2[38][17] = 4'hD;
    SS2[39][17] = 4'h0;
    SS2[40][17] = 4'h0;
    SS2[41][17] = 4'h0;
    SS2[42][17] = 4'h0;
    SS2[43][17] = 4'h0;
    SS2[44][17] = 4'h0;
    SS2[45][17] = 4'h0;
    SS2[46][17] = 4'h0;
    SS2[47][17] = 4'h0;
    SS2[0][18] = 4'h0;
    SS2[1][18] = 4'h0;
    SS2[2][18] = 4'h0;
    SS2[3][18] = 4'h0;
    SS2[4][18] = 4'h0;
    SS2[5][18] = 4'h0;
    SS2[6][18] = 4'hE;
    SS2[7][18] = 4'hE;
    SS2[8][18] = 4'hE;
    SS2[9][18] = 4'hE;
    SS2[10][18] = 4'hE;
    SS2[11][18] = 4'hE;
    SS2[12][18] = 4'hE;
    SS2[13][18] = 4'hE;
    SS2[14][18] = 4'hD;
    SS2[15][18] = 4'hD;
    SS2[16][18] = 4'hD;
    SS2[17][18] = 4'hE;
    SS2[18][18] = 4'hD;
    SS2[19][18] = 4'hD;
    SS2[20][18] = 4'hD;
    SS2[21][18] = 4'hC;
    SS2[22][18] = 4'hC;
    SS2[23][18] = 4'hD;
    SS2[24][18] = 4'hD;
    SS2[25][18] = 4'hA;
    SS2[26][18] = 4'hA;
    SS2[27][18] = 4'hC;
    SS2[28][18] = 4'hC;
    SS2[29][18] = 4'hC;
    SS2[30][18] = 4'hC;
    SS2[31][18] = 4'hC;
    SS2[32][18] = 4'hC;
    SS2[33][18] = 4'hC;
    SS2[34][18] = 4'hD;
    SS2[35][18] = 4'hD;
    SS2[36][18] = 4'hD;
    SS2[37][18] = 4'hD;
    SS2[38][18] = 4'h0;
    SS2[39][18] = 4'h0;
    SS2[40][18] = 4'h0;
    SS2[41][18] = 4'h0;
    SS2[42][18] = 4'h0;
    SS2[43][18] = 4'h0;
    SS2[44][18] = 4'h0;
    SS2[45][18] = 4'h0;
    SS2[46][18] = 4'h0;
    SS2[47][18] = 4'h0;
    SS2[0][19] = 4'h0;
    SS2[1][19] = 4'h0;
    SS2[2][19] = 4'h0;
    SS2[3][19] = 4'h0;
    SS2[4][19] = 4'h0;
    SS2[5][19] = 4'h0;
    SS2[6][19] = 4'h0;
    SS2[7][19] = 4'hE;
    SS2[8][19] = 4'hE;
    SS2[9][19] = 4'hE;
    SS2[10][19] = 4'hE;
    SS2[11][19] = 4'hE;
    SS2[12][19] = 4'hE;
    SS2[13][19] = 4'hE;
    SS2[14][19] = 4'hE;
    SS2[15][19] = 4'hD;
    SS2[16][19] = 4'hE;
    SS2[17][19] = 4'hE;
    SS2[18][19] = 4'hE;
    SS2[19][19] = 4'hD;
    SS2[20][19] = 4'hC;
    SS2[21][19] = 4'hC;
    SS2[22][19] = 4'hC;
    SS2[23][19] = 4'hC;
    SS2[24][19] = 4'hA;
    SS2[25][19] = 4'hA;
    SS2[26][19] = 4'hA;
    SS2[27][19] = 4'hA;
    SS2[28][19] = 4'hC;
    SS2[29][19] = 4'hC;
    SS2[30][19] = 4'hC;
    SS2[31][19] = 4'hC;
    SS2[32][19] = 4'hC;
    SS2[33][19] = 4'hD;
    SS2[34][19] = 4'hD;
    SS2[35][19] = 4'hD;
    SS2[36][19] = 4'hD;
    SS2[37][19] = 4'h0;
    SS2[38][19] = 4'h0;
    SS2[39][19] = 4'h0;
    SS2[40][19] = 4'h0;
    SS2[41][19] = 4'h0;
    SS2[42][19] = 4'h0;
    SS2[43][19] = 4'h0;
    SS2[44][19] = 4'h0;
    SS2[45][19] = 4'h0;
    SS2[46][19] = 4'h0;
    SS2[47][19] = 4'h0;
    SS2[0][20] = 4'h0;
    SS2[1][20] = 4'h0;
    SS2[2][20] = 4'h0;
    SS2[3][20] = 4'h0;
    SS2[4][20] = 4'h0;
    SS2[5][20] = 4'h0;
    SS2[6][20] = 4'h0;
    SS2[7][20] = 4'h0;
    SS2[8][20] = 4'hE;
    SS2[9][20] = 4'hE;
    SS2[10][20] = 4'hE;
    SS2[11][20] = 4'hC;
    SS2[12][20] = 4'hE;
    SS2[13][20] = 4'hE;
    SS2[14][20] = 4'hE;
    SS2[15][20] = 4'hC;
    SS2[16][20] = 4'hE;
    SS2[17][20] = 4'hE;
    SS2[18][20] = 4'hE;
    SS2[19][20] = 4'hC;
    SS2[20][20] = 4'hC;
    SS2[21][20] = 4'hC;
    SS2[22][20] = 4'hC;
    SS2[23][20] = 4'hD;
    SS2[24][20] = 4'hD;
    SS2[25][20] = 4'hA;
    SS2[26][20] = 4'hA;
    SS2[27][20] = 4'hA;
    SS2[28][20] = 4'hA;
    SS2[29][20] = 4'hC;
    SS2[30][20] = 4'hC;
    SS2[31][20] = 4'hC;
    SS2[32][20] = 4'hC;
    SS2[33][20] = 4'hD;
    SS2[34][20] = 4'hD;
    SS2[35][20] = 4'hD;
    SS2[36][20] = 4'h0;
    SS2[37][20] = 4'h0;
    SS2[38][20] = 4'h0;
    SS2[39][20] = 4'h0;
    SS2[40][20] = 4'h0;
    SS2[41][20] = 4'h0;
    SS2[42][20] = 4'h0;
    SS2[43][20] = 4'h0;
    SS2[44][20] = 4'h0;
    SS2[45][20] = 4'h0;
    SS2[46][20] = 4'h0;
    SS2[47][20] = 4'h0;
    SS2[0][21] = 4'h0;
    SS2[1][21] = 4'h0;
    SS2[2][21] = 4'h0;
    SS2[3][21] = 4'h0;
    SS2[4][21] = 4'h0;
    SS2[5][21] = 4'h0;
    SS2[6][21] = 4'h0;
    SS2[7][21] = 4'h0;
    SS2[8][21] = 4'h0;
    SS2[9][21] = 4'hE;
    SS2[10][21] = 4'hC;
    SS2[11][21] = 4'hC;
    SS2[12][21] = 4'hC;
    SS2[13][21] = 4'hE;
    SS2[14][21] = 4'hC;
    SS2[15][21] = 4'hC;
    SS2[16][21] = 4'hC;
    SS2[17][21] = 4'hE;
    SS2[18][21] = 4'hC;
    SS2[19][21] = 4'hC;
    SS2[20][21] = 4'hC;
    SS2[21][21] = 4'hC;
    SS2[22][21] = 4'hD;
    SS2[23][21] = 4'hD;
    SS2[24][21] = 4'hD;
    SS2[25][21] = 4'hD;
    SS2[26][21] = 4'hA;
    SS2[27][21] = 4'hA;
    SS2[28][21] = 4'hA;
    SS2[29][21] = 4'hA;
    SS2[30][21] = 4'hC;
    SS2[31][21] = 4'hC;
    SS2[32][21] = 4'hC;
    SS2[33][21] = 4'hC;
    SS2[34][21] = 4'hD;
    SS2[35][21] = 4'h0;
    SS2[36][21] = 4'h0;
    SS2[37][21] = 4'h0;
    SS2[38][21] = 4'h0;
    SS2[39][21] = 4'h0;
    SS2[40][21] = 4'h0;
    SS2[41][21] = 4'h0;
    SS2[42][21] = 4'h0;
    SS2[43][21] = 4'h0;
    SS2[44][21] = 4'h0;
    SS2[45][21] = 4'h0;
    SS2[46][21] = 4'h0;
    SS2[47][21] = 4'h0;
    SS2[0][22] = 4'h0;
    SS2[1][22] = 4'h0;
    SS2[2][22] = 4'h0;
    SS2[3][22] = 4'h0;
    SS2[4][22] = 4'h0;
    SS2[5][22] = 4'h0;
    SS2[6][22] = 4'h0;
    SS2[7][22] = 4'h0;
    SS2[8][22] = 4'hD;
    SS2[9][22] = 4'hC;
    SS2[10][22] = 4'hC;
    SS2[11][22] = 4'hC;
    SS2[12][22] = 4'hC;
    SS2[13][22] = 4'hC;
    SS2[14][22] = 4'hC;
    SS2[15][22] = 4'hC;
    SS2[16][22] = 4'hC;
    SS2[17][22] = 4'hC;
    SS2[18][22] = 4'hC;
    SS2[19][22] = 4'hC;
    SS2[20][22] = 4'hC;
    SS2[21][22] = 4'hC;
    SS2[22][22] = 4'hC;
    SS2[23][22] = 4'hD;
    SS2[24][22] = 4'hD;
    SS2[25][22] = 4'hD;
    SS2[26][22] = 4'hD;
    SS2[27][22] = 4'hA;
    SS2[28][22] = 4'hA;
    SS2[29][22] = 4'hA;
    SS2[30][22] = 4'hD;
    SS2[31][22] = 4'hC;
    SS2[32][22] = 4'hC;
    SS2[33][22] = 4'hC;
    SS2[34][22] = 4'h0;
    SS2[35][22] = 4'h0;
    SS2[36][22] = 4'h0;
    SS2[37][22] = 4'h0;
    SS2[38][22] = 4'h0;
    SS2[39][22] = 4'h0;
    SS2[40][22] = 4'h0;
    SS2[41][22] = 4'h0;
    SS2[42][22] = 4'h0;
    SS2[43][22] = 4'h0;
    SS2[44][22] = 4'h0;
    SS2[45][22] = 4'h0;
    SS2[46][22] = 4'h0;
    SS2[47][22] = 4'h0;
    SS2[0][23] = 4'h0;
    SS2[1][23] = 4'h0;
    SS2[2][23] = 4'h0;
    SS2[3][23] = 4'h0;
    SS2[4][23] = 4'h0;
    SS2[5][23] = 4'h0;
    SS2[6][23] = 4'h0;
    SS2[7][23] = 4'hD;
    SS2[8][23] = 4'hC;
    SS2[9][23] = 4'hC;
    SS2[10][23] = 4'hC;
    SS2[11][23] = 4'hC;
    SS2[12][23] = 4'hC;
    SS2[13][23] = 4'hC;
    SS2[14][23] = 4'hC;
    SS2[15][23] = 4'hC;
    SS2[16][23] = 4'hC;
    SS2[17][23] = 4'hC;
    SS2[18][23] = 4'hC;
    SS2[19][23] = 4'hC;
    SS2[20][23] = 4'hC;
    SS2[21][23] = 4'hC;
    SS2[22][23] = 4'hC;
    SS2[23][23] = 4'hC;
    SS2[24][23] = 4'hD;
    SS2[25][23] = 4'hD;
    SS2[26][23] = 4'hD;
    SS2[27][23] = 4'hD;
    SS2[28][23] = 4'hA;
    SS2[29][23] = 4'hD;
    SS2[30][23] = 4'hD;
    SS2[31][23] = 4'hD;
    SS2[32][23] = 4'hC;
    SS2[33][23] = 4'h0;
    SS2[34][23] = 4'h0;
    SS2[35][23] = 4'h0;
    SS2[36][23] = 4'h0;
    SS2[37][23] = 4'h0;
    SS2[38][23] = 4'h0;
    SS2[39][23] = 4'h0;
    SS2[40][23] = 4'h0;
    SS2[41][23] = 4'h0;
    SS2[42][23] = 4'h0;
    SS2[43][23] = 4'h0;
    SS2[44][23] = 4'h0;
    SS2[45][23] = 4'h0;
    SS2[46][23] = 4'h0;
    SS2[47][23] = 4'h0;
    SS2[0][24] = 4'h0;
    SS2[1][24] = 4'h0;
    SS2[2][24] = 4'hC;
    SS2[3][24] = 4'h0;
    SS2[4][24] = 4'h0;
    SS2[5][24] = 4'h0;
    SS2[6][24] = 4'h0;
    SS2[7][24] = 4'hC;
    SS2[8][24] = 4'hC;
    SS2[9][24] = 4'hC;
    SS2[10][24] = 4'hC;
    SS2[11][24] = 4'hC;
    SS2[12][24] = 4'hC;
    SS2[13][24] = 4'hC;
    SS2[14][24] = 4'hC;
    SS2[15][24] = 4'hC;
    SS2[16][24] = 4'hC;
    SS2[17][24] = 4'hC;
    SS2[18][24] = 4'hC;
    SS2[19][24] = 4'hD;
    SS2[20][24] = 4'hC;
    SS2[21][24] = 4'hC;
    SS2[22][24] = 4'hC;
    SS2[23][24] = 4'hC;
    SS2[24][24] = 4'hC;
    SS2[25][24] = 4'hD;
    SS2[26][24] = 4'hD;
    SS2[27][24] = 4'hD;
    SS2[28][24] = 4'hC;
    SS2[29][24] = 4'hD;
    SS2[30][24] = 4'hD;
    SS2[31][24] = 4'hD;
    SS2[32][24] = 4'hD;
    SS2[33][24] = 4'h0;
    SS2[34][24] = 4'h0;
    SS2[35][24] = 4'h0;
    SS2[36][24] = 4'h0;
    SS2[37][24] = 4'h0;
    SS2[38][24] = 4'h0;
    SS2[39][24] = 4'h0;
    SS2[40][24] = 4'h0;
    SS2[41][24] = 4'h0;
    SS2[42][24] = 4'h0;
    SS2[43][24] = 4'h0;
    SS2[44][24] = 4'h0;
    SS2[45][24] = 4'h0;
    SS2[46][24] = 4'h0;
    SS2[47][24] = 4'h0;
    SS2[0][25] = 4'h0;
    SS2[1][25] = 4'hC;
    SS2[2][25] = 4'hC;
    SS2[3][25] = 4'hC;
    SS2[4][25] = 4'h0;
    SS2[5][25] = 4'h0;
    SS2[6][25] = 4'hC;
    SS2[7][25] = 4'hC;
    SS2[8][25] = 4'hC;
    SS2[9][25] = 4'hC;
    SS2[10][25] = 4'hC;
    SS2[11][25] = 4'hC;
    SS2[12][25] = 4'hC;
    SS2[13][25] = 4'hC;
    SS2[14][25] = 4'hC;
    SS2[15][25] = 4'hC;
    SS2[16][25] = 4'hC;
    SS2[17][25] = 4'hC;
    SS2[18][25] = 4'hD;
    SS2[19][25] = 4'hD;
    SS2[20][25] = 4'hD;
    SS2[21][25] = 4'hC;
    SS2[22][25] = 4'hC;
    SS2[23][25] = 4'hC;
    SS2[24][25] = 4'hC;
    SS2[25][25] = 4'hC;
    SS2[26][25] = 4'hD;
    SS2[27][25] = 4'hC;
    SS2[28][25] = 4'hC;
    SS2[29][25] = 4'hC;
    SS2[30][25] = 4'hD;
    SS2[31][25] = 4'hD;
    SS2[32][25] = 4'hD;
    SS2[33][25] = 4'hD;
    SS2[34][25] = 4'h0;
    SS2[35][25] = 4'h0;
    SS2[36][25] = 4'h0;
    SS2[37][25] = 4'h0;
    SS2[38][25] = 4'h0;
    SS2[39][25] = 4'h0;
    SS2[40][25] = 4'h0;
    SS2[41][25] = 4'h0;
    SS2[42][25] = 4'h0;
    SS2[43][25] = 4'h0;
    SS2[44][25] = 4'h0;
    SS2[45][25] = 4'h0;
    SS2[46][25] = 4'h0;
    SS2[47][25] = 4'h0;
    SS2[0][26] = 4'hC;
    SS2[1][26] = 4'hC;
    SS2[2][26] = 4'hC;
    SS2[3][26] = 4'hC;
    SS2[4][26] = 4'hC;
    SS2[5][26] = 4'hC;
    SS2[6][26] = 4'hC;
    SS2[7][26] = 4'hC;
    SS2[8][26] = 4'hC;
    SS2[9][26] = 4'hD;
    SS2[10][26] = 4'hC;
    SS2[11][26] = 4'hC;
    SS2[12][26] = 4'hC;
    SS2[13][26] = 4'hD;
    SS2[14][26] = 4'hC;
    SS2[15][26] = 4'hC;
    SS2[16][26] = 4'hC;
    SS2[17][26] = 4'hE;
    SS2[18][26] = 4'hD;
    SS2[19][26] = 4'hD;
    SS2[20][26] = 4'hD;
    SS2[21][26] = 4'hD;
    SS2[22][26] = 4'hC;
    SS2[23][26] = 4'hC;
    SS2[24][26] = 4'hC;
    SS2[25][26] = 4'hC;
    SS2[26][26] = 4'hC;
    SS2[27][26] = 4'hC;
    SS2[28][26] = 4'hC;
    SS2[29][26] = 4'hC;
    SS2[30][26] = 4'hD;
    SS2[31][26] = 4'hD;
    SS2[32][26] = 4'hD;
    SS2[33][26] = 4'hD;
    SS2[34][26] = 4'h3;
    SS2[35][26] = 4'h0;
    SS2[36][26] = 4'h0;
    SS2[37][26] = 4'h0;
    SS2[38][26] = 4'h0;
    SS2[39][26] = 4'h0;
    SS2[40][26] = 4'h0;
    SS2[41][26] = 4'h0;
    SS2[42][26] = 4'h0;
    SS2[43][26] = 4'h0;
    SS2[44][26] = 4'h0;
    SS2[45][26] = 4'h0;
    SS2[46][26] = 4'h0;
    SS2[47][26] = 4'h0;
    SS2[0][27] = 4'hC;
    SS2[1][27] = 4'hC;
    SS2[2][27] = 4'hC;
    SS2[3][27] = 4'hC;
    SS2[4][27] = 4'hC;
    SS2[5][27] = 4'hC;
    SS2[6][27] = 4'hC;
    SS2[7][27] = 4'hC;
    SS2[8][27] = 4'hD;
    SS2[9][27] = 4'hD;
    SS2[10][27] = 4'hD;
    SS2[11][27] = 4'hC;
    SS2[12][27] = 4'hD;
    SS2[13][27] = 4'hD;
    SS2[14][27] = 4'hD;
    SS2[15][27] = 4'hC;
    SS2[16][27] = 4'hE;
    SS2[17][27] = 4'hE;
    SS2[18][27] = 4'hE;
    SS2[19][27] = 4'hD;
    SS2[20][27] = 4'hD;
    SS2[21][27] = 4'hD;
    SS2[22][27] = 4'hD;
    SS2[23][27] = 4'hC;
    SS2[24][27] = 4'hC;
    SS2[25][27] = 4'hC;
    SS2[26][27] = 4'hC;
    SS2[27][27] = 4'hC;
    SS2[28][27] = 4'hC;
    SS2[29][27] = 4'hD;
    SS2[30][27] = 4'hD;
    SS2[31][27] = 4'hD;
    SS2[32][27] = 4'hD;
    SS2[33][27] = 4'h3;
    SS2[34][27] = 4'h3;
    SS2[35][27] = 4'h3;
    SS2[36][27] = 4'h0;
    SS2[37][27] = 4'h0;
    SS2[38][27] = 4'h0;
    SS2[39][27] = 4'h0;
    SS2[40][27] = 4'h0;
    SS2[41][27] = 4'h0;
    SS2[42][27] = 4'h0;
    SS2[43][27] = 4'h0;
    SS2[44][27] = 4'h0;
    SS2[45][27] = 4'h0;
    SS2[46][27] = 4'h0;
    SS2[47][27] = 4'h0;
    SS2[0][28] = 4'hC;
    SS2[1][28] = 4'hC;
    SS2[2][28] = 4'hC;
    SS2[3][28] = 4'hC;
    SS2[4][28] = 4'hC;
    SS2[5][28] = 4'hC;
    SS2[6][28] = 4'hC;
    SS2[7][28] = 4'hD;
    SS2[8][28] = 4'hD;
    SS2[9][28] = 4'hD;
    SS2[10][28] = 4'hD;
    SS2[11][28] = 4'hD;
    SS2[12][28] = 4'hD;
    SS2[13][28] = 4'hD;
    SS2[14][28] = 4'hD;
    SS2[15][28] = 4'hE;
    SS2[16][28] = 4'hE;
    SS2[17][28] = 4'hE;
    SS2[18][28] = 4'hE;
    SS2[19][28] = 4'hE;
    SS2[20][28] = 4'hD;
    SS2[21][28] = 4'hD;
    SS2[22][28] = 4'hD;
    SS2[23][28] = 4'hD;
    SS2[24][28] = 4'hC;
    SS2[25][28] = 4'hC;
    SS2[26][28] = 4'hC;
    SS2[27][28] = 4'hC;
    SS2[28][28] = 4'hD;
    SS2[29][28] = 4'hD;
    SS2[30][28] = 4'hD;
    SS2[31][28] = 4'hD;
    SS2[32][28] = 4'hD;
    SS2[33][28] = 4'h3;
    SS2[34][28] = 4'h3;
    SS2[35][28] = 4'h3;
    SS2[36][28] = 4'h2;
    SS2[37][28] = 4'h0;
    SS2[38][28] = 4'h0;
    SS2[39][28] = 4'h0;
    SS2[40][28] = 4'h0;
    SS2[41][28] = 4'h0;
    SS2[42][28] = 4'h0;
    SS2[43][28] = 4'h0;
    SS2[44][28] = 4'h0;
    SS2[45][28] = 4'h0;
    SS2[46][28] = 4'h0;
    SS2[47][28] = 4'h0;
    SS2[0][29] = 4'hC;
    SS2[1][29] = 4'hC;
    SS2[2][29] = 4'hD;
    SS2[3][29] = 4'hD;
    SS2[4][29] = 4'hC;
    SS2[5][29] = 4'hC;
    SS2[6][29] = 4'hE;
    SS2[7][29] = 4'hE;
    SS2[8][29] = 4'hD;
    SS2[9][29] = 4'hD;
    SS2[10][29] = 4'hE;
    SS2[11][29] = 4'hE;
    SS2[12][29] = 4'hD;
    SS2[13][29] = 4'hD;
    SS2[14][29] = 4'hE;
    SS2[15][29] = 4'hE;
    SS2[16][29] = 4'hE;
    SS2[17][29] = 4'hE;
    SS2[18][29] = 4'hE;
    SS2[19][29] = 4'hE;
    SS2[20][29] = 4'hE;
    SS2[21][29] = 4'hD;
    SS2[22][29] = 4'hD;
    SS2[23][29] = 4'hC;
    SS2[24][29] = 4'hC;
    SS2[25][29] = 4'hC;
    SS2[26][29] = 4'hC;
    SS2[27][29] = 4'hE;
    SS2[28][29] = 4'hE;
    SS2[29][29] = 4'hD;
    SS2[30][29] = 4'hD;
    SS2[31][29] = 4'hD;
    SS2[32][29] = 4'hD;
    SS2[33][29] = 4'hD;
    SS2[34][29] = 4'h3;
    SS2[35][29] = 4'h2;
    SS2[36][29] = 4'h0;
    SS2[37][29] = 4'h0;
    SS2[38][29] = 4'h0;
    SS2[39][29] = 4'h0;
    SS2[40][29] = 4'h0;
    SS2[41][29] = 4'h0;
    SS2[42][29] = 4'h0;
    SS2[43][29] = 4'h0;
    SS2[44][29] = 4'h0;
    SS2[45][29] = 4'h0;
    SS2[46][29] = 4'h0;
    SS2[47][29] = 4'h0;
    SS2[0][30] = 4'hE;
    SS2[1][30] = 4'hD;
    SS2[2][30] = 4'hD;
    SS2[3][30] = 4'hD;
    SS2[4][30] = 4'hD;
    SS2[5][30] = 4'hE;
    SS2[6][30] = 4'hE;
    SS2[7][30] = 4'hE;
    SS2[8][30] = 4'hE;
    SS2[9][30] = 4'hE;
    SS2[10][30] = 4'hE;
    SS2[11][30] = 4'hE;
    SS2[12][30] = 4'hE;
    SS2[13][30] = 4'h0;
    SS2[14][30] = 4'hE;
    SS2[15][30] = 4'hE;
    SS2[16][30] = 4'hE;
    SS2[17][30] = 4'hE;
    SS2[18][30] = 4'hE;
    SS2[19][30] = 4'hE;
    SS2[20][30] = 4'hE;
    SS2[21][30] = 4'hE;
    SS2[22][30] = 4'hC;
    SS2[23][30] = 4'hC;
    SS2[24][30] = 4'hC;
    SS2[25][30] = 4'hC;
    SS2[26][30] = 4'hE;
    SS2[27][30] = 4'hE;
    SS2[28][30] = 4'hE;
    SS2[29][30] = 4'hE;
    SS2[30][30] = 4'hD;
    SS2[31][30] = 4'hD;
    SS2[32][30] = 4'hD;
    SS2[33][30] = 4'hD;
    SS2[34][30] = 4'h0;
    SS2[35][30] = 4'h0;
    SS2[36][30] = 4'h0;
    SS2[37][30] = 4'h0;
    SS2[38][30] = 4'h0;
    SS2[39][30] = 4'h0;
    SS2[40][30] = 4'h0;
    SS2[41][30] = 4'h0;
    SS2[42][30] = 4'h0;
    SS2[43][30] = 4'h0;
    SS2[44][30] = 4'h0;
    SS2[45][30] = 4'h0;
    SS2[46][30] = 4'h0;
    SS2[47][30] = 4'h0;
    SS2[0][31] = 4'h0;
    SS2[1][31] = 4'h0;
    SS2[2][31] = 4'hD;
    SS2[3][31] = 4'hD;
    SS2[4][31] = 4'h0;
    SS2[5][31] = 4'h0;
    SS2[6][31] = 4'hE;
    SS2[7][31] = 4'hE;
    SS2[8][31] = 4'h0;
    SS2[9][31] = 4'h0;
    SS2[10][31] = 4'hE;
    SS2[11][31] = 4'hE;
    SS2[12][31] = 4'h0;
    SS2[13][31] = 4'h0;
    SS2[14][31] = 4'h0;
    SS2[15][31] = 4'hE;
    SS2[16][31] = 4'hE;
    SS2[17][31] = 4'hE;
    SS2[18][31] = 4'hE;
    SS2[19][31] = 4'hE;
    SS2[20][31] = 4'hE;
    SS2[21][31] = 4'hC;
    SS2[22][31] = 4'hC;
    SS2[23][31] = 4'hC;
    SS2[24][31] = 4'hC;
    SS2[25][31] = 4'hC;
    SS2[26][31] = 4'hC;
    SS2[27][31] = 4'hE;
    SS2[28][31] = 4'hE;
    SS2[29][31] = 4'hD;
    SS2[30][31] = 4'hD;
    SS2[31][31] = 4'hD;
    SS2[32][31] = 4'hD;
    SS2[33][31] = 4'h0;
    SS2[34][31] = 4'h0;
    SS2[35][31] = 4'h0;
    SS2[36][31] = 4'h0;
    SS2[37][31] = 4'h0;
    SS2[38][31] = 4'h0;
    SS2[39][31] = 4'h0;
    SS2[40][31] = 4'h0;
    SS2[41][31] = 4'h0;
    SS2[42][31] = 4'h0;
    SS2[43][31] = 4'h0;
    SS2[44][31] = 4'h0;
    SS2[45][31] = 4'h0;
    SS2[46][31] = 4'h0;
    SS2[47][31] = 4'h0;
    SS2[0][32] = 4'h0;
    SS2[1][32] = 4'h0;
    SS2[2][32] = 4'h0;
    SS2[3][32] = 4'h0;
    SS2[4][32] = 4'h0;
    SS2[5][32] = 4'h0;
    SS2[6][32] = 4'h0;
    SS2[7][32] = 4'h0;
    SS2[8][32] = 4'h0;
    SS2[9][32] = 4'h0;
    SS2[10][32] = 4'h0;
    SS2[11][32] = 4'h0;
    SS2[12][32] = 4'h0;
    SS2[13][32] = 4'h0;
    SS2[14][32] = 4'h0;
    SS2[15][32] = 4'hF;
    SS2[16][32] = 4'hE;
    SS2[17][32] = 4'hE;
    SS2[18][32] = 4'hE;
    SS2[19][32] = 4'hE;
    SS2[20][32] = 4'hC;
    SS2[21][32] = 4'hC;
    SS2[22][32] = 4'hC;
    SS2[23][32] = 4'hC;
    SS2[24][32] = 4'hC;
    SS2[25][32] = 4'hC;
    SS2[26][32] = 4'hC;
    SS2[27][32] = 4'hC;
    SS2[28][32] = 4'hD;
    SS2[29][32] = 4'hD;
    SS2[30][32] = 4'hD;
    SS2[31][32] = 4'hD;
    SS2[32][32] = 4'hD;
    SS2[33][32] = 4'h0;
    SS2[34][32] = 4'h0;
    SS2[35][32] = 4'h0;
    SS2[36][32] = 4'h0;
    SS2[37][32] = 4'h0;
    SS2[38][32] = 4'h0;
    SS2[39][32] = 4'h0;
    SS2[40][32] = 4'h0;
    SS2[41][32] = 4'h0;
    SS2[42][32] = 4'h0;
    SS2[43][32] = 4'h0;
    SS2[44][32] = 4'h0;
    SS2[45][32] = 4'h0;
    SS2[46][32] = 4'h0;
    SS2[47][32] = 4'h0;
    SS2[0][33] = 4'h0;
    SS2[1][33] = 4'h0;
    SS2[2][33] = 4'h0;
    SS2[3][33] = 4'h0;
    SS2[4][33] = 4'h0;
    SS2[5][33] = 4'h0;
    SS2[6][33] = 4'h0;
    SS2[7][33] = 4'h0;
    SS2[8][33] = 4'h0;
    SS2[9][33] = 4'h0;
    SS2[10][33] = 4'h0;
    SS2[11][33] = 4'h0;
    SS2[12][33] = 4'h0;
    SS2[13][33] = 4'h0;
    SS2[14][33] = 4'h0;
    SS2[15][33] = 4'h0;
    SS2[16][33] = 4'h0;
    SS2[17][33] = 4'hE;
    SS2[18][33] = 4'hE;
    SS2[19][33] = 4'hD;
    SS2[20][33] = 4'hD;
    SS2[21][33] = 4'hC;
    SS2[22][33] = 4'hC;
    SS2[23][33] = 4'hC;
    SS2[24][33] = 4'hC;
    SS2[25][33] = 4'hC;
    SS2[26][33] = 4'hC;
    SS2[27][33] = 4'hE;
    SS2[28][33] = 4'hE;
    SS2[29][33] = 4'hD;
    SS2[30][33] = 4'hD;
    SS2[31][33] = 4'hD;
    SS2[32][33] = 4'hD;
    SS2[33][33] = 4'hE;
    SS2[34][33] = 4'h0;
    SS2[35][33] = 4'h0;
    SS2[36][33] = 4'h0;
    SS2[37][33] = 4'h0;
    SS2[38][33] = 4'h0;
    SS2[39][33] = 4'h0;
    SS2[40][33] = 4'h0;
    SS2[41][33] = 4'h0;
    SS2[42][33] = 4'h0;
    SS2[43][33] = 4'h0;
    SS2[44][33] = 4'h0;
    SS2[45][33] = 4'h0;
    SS2[46][33] = 4'h0;
    SS2[47][33] = 4'h0;
    SS2[0][34] = 4'h0;
    SS2[1][34] = 4'h0;
    SS2[2][34] = 4'h0;
    SS2[3][34] = 4'h0;
    SS2[4][34] = 4'h0;
    SS2[5][34] = 4'h0;
    SS2[6][34] = 4'h0;
    SS2[7][34] = 4'h0;
    SS2[8][34] = 4'h0;
    SS2[9][34] = 4'h0;
    SS2[10][34] = 4'h0;
    SS2[11][34] = 4'h0;
    SS2[12][34] = 4'h0;
    SS2[13][34] = 4'h0;
    SS2[14][34] = 4'h0;
    SS2[15][34] = 4'h0;
    SS2[16][34] = 4'h0;
    SS2[17][34] = 4'h0;
    SS2[18][34] = 4'hD;
    SS2[19][34] = 4'hD;
    SS2[20][34] = 4'hD;
    SS2[21][34] = 4'hD;
    SS2[22][34] = 4'hC;
    SS2[23][34] = 4'hC;
    SS2[24][34] = 4'hC;
    SS2[25][34] = 4'hC;
    SS2[26][34] = 4'hE;
    SS2[27][34] = 4'hE;
    SS2[28][34] = 4'hE;
    SS2[29][34] = 4'hE;
    SS2[30][34] = 4'hD;
    SS2[31][34] = 4'hD;
    SS2[32][34] = 4'hD;
    SS2[33][34] = 4'hD;
    SS2[34][34] = 4'hE;
    SS2[35][34] = 4'h0;
    SS2[36][34] = 4'h0;
    SS2[37][34] = 4'h0;
    SS2[38][34] = 4'h0;
    SS2[39][34] = 4'h0;
    SS2[40][34] = 4'h0;
    SS2[41][34] = 4'h0;
    SS2[42][34] = 4'h0;
    SS2[43][34] = 4'h0;
    SS2[44][34] = 4'h0;
    SS2[45][34] = 4'h0;
    SS2[46][34] = 4'h0;
    SS2[47][34] = 4'h0;
    SS2[0][35] = 4'h0;
    SS2[1][35] = 4'h0;
    SS2[2][35] = 4'h0;
    SS2[3][35] = 4'h0;
    SS2[4][35] = 4'h0;
    SS2[5][35] = 4'h0;
    SS2[6][35] = 4'h0;
    SS2[7][35] = 4'h0;
    SS2[8][35] = 4'h0;
    SS2[9][35] = 4'h0;
    SS2[10][35] = 4'h0;
    SS2[11][35] = 4'h0;
    SS2[12][35] = 4'h0;
    SS2[13][35] = 4'h0;
    SS2[14][35] = 4'h0;
    SS2[15][35] = 4'h0;
    SS2[16][35] = 4'h0;
    SS2[17][35] = 4'hE;
    SS2[18][35] = 4'hD;
    SS2[19][35] = 4'hD;
    SS2[20][35] = 4'hD;
    SS2[21][35] = 4'hC;
    SS2[22][35] = 4'hC;
    SS2[23][35] = 4'hC;
    SS2[24][35] = 4'hC;
    SS2[25][35] = 4'hC;
    SS2[26][35] = 4'hC;
    SS2[27][35] = 4'hE;
    SS2[28][35] = 4'hE;
    SS2[29][35] = 4'hE;
    SS2[30][35] = 4'hE;
    SS2[31][35] = 4'hD;
    SS2[32][35] = 4'hD;
    SS2[33][35] = 4'hD;
    SS2[34][35] = 4'h3;
    SS2[35][35] = 4'h2;
    SS2[36][35] = 4'h0;
    SS2[37][35] = 4'h0;
    SS2[38][35] = 4'h0;
    SS2[39][35] = 4'h0;
    SS2[40][35] = 4'h0;
    SS2[41][35] = 4'h0;
    SS2[42][35] = 4'h0;
    SS2[43][35] = 4'h0;
    SS2[44][35] = 4'h0;
    SS2[45][35] = 4'h0;
    SS2[46][35] = 4'h0;
    SS2[47][35] = 4'h0;
    SS2[0][36] = 4'h0;
    SS2[1][36] = 4'h0;
    SS2[2][36] = 4'h0;
    SS2[3][36] = 4'h0;
    SS2[4][36] = 4'h0;
    SS2[5][36] = 4'h0;
    SS2[6][36] = 4'h0;
    SS2[7][36] = 4'h0;
    SS2[8][36] = 4'h0;
    SS2[9][36] = 4'h0;
    SS2[10][36] = 4'h0;
    SS2[11][36] = 4'h0;
    SS2[12][36] = 4'h0;
    SS2[13][36] = 4'h0;
    SS2[14][36] = 4'h0;
    SS2[15][36] = 4'h0;
    SS2[16][36] = 4'hE;
    SS2[17][36] = 4'hE;
    SS2[18][36] = 4'hE;
    SS2[19][36] = 4'hD;
    SS2[20][36] = 4'hC;
    SS2[21][36] = 4'hC;
    SS2[22][36] = 4'hC;
    SS2[23][36] = 4'hC;
    SS2[24][36] = 4'hC;
    SS2[25][36] = 4'hC;
    SS2[26][36] = 4'hC;
    SS2[27][36] = 4'hC;
    SS2[28][36] = 4'hE;
    SS2[29][36] = 4'hE;
    SS2[30][36] = 4'hE;
    SS2[31][36] = 4'hE;
    SS2[32][36] = 4'hD;
    SS2[33][36] = 4'h3;
    SS2[34][36] = 4'h3;
    SS2[35][36] = 4'h3;
    SS2[36][36] = 4'h2;
    SS2[37][36] = 4'h0;
    SS2[38][36] = 4'h0;
    SS2[39][36] = 4'h0;
    SS2[40][36] = 4'h0;
    SS2[41][36] = 4'h0;
    SS2[42][36] = 4'h0;
    SS2[43][36] = 4'h0;
    SS2[44][36] = 4'h0;
    SS2[45][36] = 4'h0;
    SS2[46][36] = 4'h0;
    SS2[47][36] = 4'h0;
    SS2[0][37] = 4'h0;
    SS2[1][37] = 4'h0;
    SS2[2][37] = 4'h0;
    SS2[3][37] = 4'h0;
    SS2[4][37] = 4'h0;
    SS2[5][37] = 4'h0;
    SS2[6][37] = 4'h0;
    SS2[7][37] = 4'h0;
    SS2[8][37] = 4'h0;
    SS2[9][37] = 4'h0;
    SS2[10][37] = 4'h0;
    SS2[11][37] = 4'h0;
    SS2[12][37] = 4'h0;
    SS2[13][37] = 4'h0;
    SS2[14][37] = 4'h0;
    SS2[15][37] = 4'h0;
    SS2[16][37] = 4'hE;
    SS2[17][37] = 4'hE;
    SS2[18][37] = 4'hE;
    SS2[19][37] = 4'hD;
    SS2[20][37] = 4'hD;
    SS2[21][37] = 4'hC;
    SS2[22][37] = 4'hC;
    SS2[23][37] = 4'hC;
    SS2[24][37] = 4'hC;
    SS2[25][37] = 4'hC;
    SS2[26][37] = 4'hC;
    SS2[27][37] = 4'hE;
    SS2[28][37] = 4'hE;
    SS2[29][37] = 4'hE;
    SS2[30][37] = 4'hE;
    SS2[31][37] = 4'hE;
    SS2[32][37] = 4'hD;
    SS2[33][37] = 4'h3;
    SS2[34][37] = 4'h3;
    SS2[35][37] = 4'h3;
    SS2[36][37] = 4'h0;
    SS2[37][37] = 4'h0;
    SS2[38][37] = 4'h0;
    SS2[39][37] = 4'h0;
    SS2[40][37] = 4'h0;
    SS2[41][37] = 4'h0;
    SS2[42][37] = 4'h0;
    SS2[43][37] = 4'h0;
    SS2[44][37] = 4'h0;
    SS2[45][37] = 4'h0;
    SS2[46][37] = 4'h0;
    SS2[47][37] = 4'h0;
    SS2[0][38] = 4'h0;
    SS2[1][38] = 4'h0;
    SS2[2][38] = 4'h0;
    SS2[3][38] = 4'h0;
    SS2[4][38] = 4'h0;
    SS2[5][38] = 4'h0;
    SS2[6][38] = 4'h0;
    SS2[7][38] = 4'h0;
    SS2[8][38] = 4'h0;
    SS2[9][38] = 4'h0;
    SS2[10][38] = 4'h0;
    SS2[11][38] = 4'h0;
    SS2[12][38] = 4'h0;
    SS2[13][38] = 4'h0;
    SS2[14][38] = 4'h0;
    SS2[15][38] = 4'h0;
    SS2[16][38] = 4'h0;
    SS2[17][38] = 4'hE;
    SS2[18][38] = 4'hD;
    SS2[19][38] = 4'hD;
    SS2[20][38] = 4'hD;
    SS2[21][38] = 4'hD;
    SS2[22][38] = 4'hC;
    SS2[23][38] = 4'hC;
    SS2[24][38] = 4'hC;
    SS2[25][38] = 4'hC;
    SS2[26][38] = 4'hE;
    SS2[27][38] = 4'hE;
    SS2[28][38] = 4'hE;
    SS2[29][38] = 4'hE;
    SS2[30][38] = 4'hE;
    SS2[31][38] = 4'hD;
    SS2[32][38] = 4'hD;
    SS2[33][38] = 4'hD;
    SS2[34][38] = 4'h3;
    SS2[35][38] = 4'h0;
    SS2[36][38] = 4'h0;
    SS2[37][38] = 4'h0;
    SS2[38][38] = 4'h0;
    SS2[39][38] = 4'h0;
    SS2[40][38] = 4'h0;
    SS2[41][38] = 4'h0;
    SS2[42][38] = 4'h0;
    SS2[43][38] = 4'h0;
    SS2[44][38] = 4'h0;
    SS2[45][38] = 4'h0;
    SS2[46][38] = 4'h0;
    SS2[47][38] = 4'h0;
    SS2[0][39] = 4'h0;
    SS2[1][39] = 4'h0;
    SS2[2][39] = 4'h0;
    SS2[3][39] = 4'h0;
    SS2[4][39] = 4'h0;
    SS2[5][39] = 4'h0;
    SS2[6][39] = 4'h0;
    SS2[7][39] = 4'h0;
    SS2[8][39] = 4'h0;
    SS2[9][39] = 4'h0;
    SS2[10][39] = 4'h0;
    SS2[11][39] = 4'h0;
    SS2[12][39] = 4'h0;
    SS2[13][39] = 4'h0;
    SS2[14][39] = 4'h0;
    SS2[15][39] = 4'h0;
    SS2[16][39] = 4'h0;
    SS2[17][39] = 4'hE;
    SS2[18][39] = 4'hD;
    SS2[19][39] = 4'hD;
    SS2[20][39] = 4'hD;
    SS2[21][39] = 4'hC;
    SS2[22][39] = 4'hC;
    SS2[23][39] = 4'hC;
    SS2[24][39] = 4'hC;
    SS2[25][39] = 4'hD;
    SS2[26][39] = 4'h0;
    SS2[27][39] = 4'hE;
    SS2[28][39] = 4'hE;
    SS2[29][39] = 4'hE;
    SS2[30][39] = 4'hE;
    SS2[31][39] = 4'hD;
    SS2[32][39] = 4'hD;
    SS2[33][39] = 4'hD;
    SS2[34][39] = 4'hD;
    SS2[35][39] = 4'h0;
    SS2[36][39] = 4'h0;
    SS2[37][39] = 4'h0;
    SS2[38][39] = 4'h0;
    SS2[39][39] = 4'h0;
    SS2[40][39] = 4'h0;
    SS2[41][39] = 4'h0;
    SS2[42][39] = 4'h0;
    SS2[43][39] = 4'h0;
    SS2[44][39] = 4'h0;
    SS2[45][39] = 4'h0;
    SS2[46][39] = 4'h0;
    SS2[47][39] = 4'h0;
    SS2[0][40] = 4'h0;
    SS2[1][40] = 4'h0;
    SS2[2][40] = 4'h0;
    SS2[3][40] = 4'h0;
    SS2[4][40] = 4'h0;
    SS2[5][40] = 4'h0;
    SS2[6][40] = 4'h0;
    SS2[7][40] = 4'h0;
    SS2[8][40] = 4'h0;
    SS2[9][40] = 4'h0;
    SS2[10][40] = 4'h0;
    SS2[11][40] = 4'h0;
    SS2[12][40] = 4'h0;
    SS2[13][40] = 4'h0;
    SS2[14][40] = 4'h0;
    SS2[15][40] = 4'h0;
    SS2[16][40] = 4'hE;
    SS2[17][40] = 4'hE;
    SS2[18][40] = 4'hE;
    SS2[19][40] = 4'hD;
    SS2[20][40] = 4'hC;
    SS2[21][40] = 4'hC;
    SS2[22][40] = 4'hC;
    SS2[23][40] = 4'hC;
    SS2[24][40] = 4'hD;
    SS2[25][40] = 4'h0;
    SS2[26][40] = 4'h0;
    SS2[27][40] = 4'h0;
    SS2[28][40] = 4'hE;
    SS2[29][40] = 4'hE;
    SS2[30][40] = 4'hE;
    SS2[31][40] = 4'hE;
    SS2[32][40] = 4'hD;
    SS2[33][40] = 4'hD;
    SS2[34][40] = 4'hD;
    SS2[35][40] = 4'hD;
    SS2[36][40] = 4'h0;
    SS2[37][40] = 4'h0;
    SS2[38][40] = 4'h0;
    SS2[39][40] = 4'h0;
    SS2[40][40] = 4'h0;
    SS2[41][40] = 4'h0;
    SS2[42][40] = 4'h0;
    SS2[43][40] = 4'h0;
    SS2[44][40] = 4'h0;
    SS2[45][40] = 4'h0;
    SS2[46][40] = 4'h0;
    SS2[47][40] = 4'h0;
    SS2[0][41] = 4'h0;
    SS2[1][41] = 4'h0;
    SS2[2][41] = 4'h0;
    SS2[3][41] = 4'h0;
    SS2[4][41] = 4'h0;
    SS2[5][41] = 4'h0;
    SS2[6][41] = 4'h0;
    SS2[7][41] = 4'h0;
    SS2[8][41] = 4'h0;
    SS2[9][41] = 4'h0;
    SS2[10][41] = 4'h0;
    SS2[11][41] = 4'h0;
    SS2[12][41] = 4'h0;
    SS2[13][41] = 4'h0;
    SS2[14][41] = 4'h0;
    SS2[15][41] = 4'h0;
    SS2[16][41] = 4'hE;
    SS2[17][41] = 4'hE;
    SS2[18][41] = 4'hE;
    SS2[19][41] = 4'hC;
    SS2[20][41] = 4'hC;
    SS2[21][41] = 4'hC;
    SS2[22][41] = 4'hC;
    SS2[23][41] = 4'h0;
    SS2[24][41] = 4'h0;
    SS2[25][41] = 4'h0;
    SS2[26][41] = 4'h0;
    SS2[27][41] = 4'h0;
    SS2[28][41] = 4'h0;
    SS2[29][41] = 4'hE;
    SS2[30][41] = 4'hE;
    SS2[31][41] = 4'hE;
    SS2[32][41] = 4'hD;
    SS2[33][41] = 4'hD;
    SS2[34][41] = 4'hD;
    SS2[35][41] = 4'hD;
    SS2[36][41] = 4'h0;
    SS2[37][41] = 4'h0;
    SS2[38][41] = 4'h0;
    SS2[39][41] = 4'h0;
    SS2[40][41] = 4'h0;
    SS2[41][41] = 4'h0;
    SS2[42][41] = 4'h0;
    SS2[43][41] = 4'h0;
    SS2[44][41] = 4'h0;
    SS2[45][41] = 4'h0;
    SS2[46][41] = 4'h0;
    SS2[47][41] = 4'h0;
    SS2[0][42] = 4'h0;
    SS2[1][42] = 4'h0;
    SS2[2][42] = 4'h0;
    SS2[3][42] = 4'h0;
    SS2[4][42] = 4'h0;
    SS2[5][42] = 4'h0;
    SS2[6][42] = 4'h0;
    SS2[7][42] = 4'h0;
    SS2[8][42] = 4'h0;
    SS2[9][42] = 4'h0;
    SS2[10][42] = 4'h0;
    SS2[11][42] = 4'h0;
    SS2[12][42] = 4'h0;
    SS2[13][42] = 4'h0;
    SS2[14][42] = 4'h0;
    SS2[15][42] = 4'h0;
    SS2[16][42] = 4'h0;
    SS2[17][42] = 4'hE;
    SS2[18][42] = 4'hC;
    SS2[19][42] = 4'hC;
    SS2[20][42] = 4'hC;
    SS2[21][42] = 4'hC;
    SS2[22][42] = 4'h0;
    SS2[23][42] = 4'h0;
    SS2[24][42] = 4'h0;
    SS2[25][42] = 4'h0;
    SS2[26][42] = 4'h0;
    SS2[27][42] = 4'h0;
    SS2[28][42] = 4'h0;
    SS2[29][42] = 4'h0;
    SS2[30][42] = 4'hE;
    SS2[31][42] = 4'hD;
    SS2[32][42] = 4'hD;
    SS2[33][42] = 4'hD;
    SS2[34][42] = 4'hD;
    SS2[35][42] = 4'h0;
    SS2[36][42] = 4'h0;
    SS2[37][42] = 4'h0;
    SS2[38][42] = 4'h0;
    SS2[39][42] = 4'h0;
    SS2[40][42] = 4'h0;
    SS2[41][42] = 4'h0;
    SS2[42][42] = 4'h0;
    SS2[43][42] = 4'h0;
    SS2[44][42] = 4'h0;
    SS2[45][42] = 4'h0;
    SS2[46][42] = 4'h0;
    SS2[47][42] = 4'h0;
    SS2[0][43] = 4'h0;
    SS2[1][43] = 4'h0;
    SS2[2][43] = 4'h0;
    SS2[3][43] = 4'h0;
    SS2[4][43] = 4'h0;
    SS2[5][43] = 4'h0;
    SS2[6][43] = 4'h0;
    SS2[7][43] = 4'h0;
    SS2[8][43] = 4'h0;
    SS2[9][43] = 4'h0;
    SS2[10][43] = 4'h0;
    SS2[11][43] = 4'h0;
    SS2[12][43] = 4'h0;
    SS2[13][43] = 4'h0;
    SS2[14][43] = 4'h0;
    SS2[15][43] = 4'h0;
    SS2[16][43] = 4'h0;
    SS2[17][43] = 4'hD;
    SS2[18][43] = 4'hC;
    SS2[19][43] = 4'hC;
    SS2[20][43] = 4'hC;
    SS2[21][43] = 4'hC;
    SS2[22][43] = 4'h0;
    SS2[23][43] = 4'h0;
    SS2[24][43] = 4'h0;
    SS2[25][43] = 4'h0;
    SS2[26][43] = 4'h0;
    SS2[27][43] = 4'h0;
    SS2[28][43] = 4'h0;
    SS2[29][43] = 4'h0;
    SS2[30][43] = 4'h0;
    SS2[31][43] = 4'hD;
    SS2[32][43] = 4'hD;
    SS2[33][43] = 4'hD;
    SS2[34][43] = 4'hD;
    SS2[35][43] = 4'h0;
    SS2[36][43] = 4'h0;
    SS2[37][43] = 4'h0;
    SS2[38][43] = 4'h0;
    SS2[39][43] = 4'h0;
    SS2[40][43] = 4'h0;
    SS2[41][43] = 4'h0;
    SS2[42][43] = 4'h0;
    SS2[43][43] = 4'h0;
    SS2[44][43] = 4'h0;
    SS2[45][43] = 4'h0;
    SS2[46][43] = 4'h0;
    SS2[47][43] = 4'h0;
    SS2[0][44] = 4'h0;
    SS2[1][44] = 4'h0;
    SS2[2][44] = 4'h0;
    SS2[3][44] = 4'h0;
    SS2[4][44] = 4'h0;
    SS2[5][44] = 4'h0;
    SS2[6][44] = 4'h0;
    SS2[7][44] = 4'h0;
    SS2[8][44] = 4'h0;
    SS2[9][44] = 4'h0;
    SS2[10][44] = 4'h0;
    SS2[11][44] = 4'h0;
    SS2[12][44] = 4'h0;
    SS2[13][44] = 4'h0;
    SS2[14][44] = 4'h0;
    SS2[15][44] = 4'h0;
    SS2[16][44] = 4'hD;
    SS2[17][44] = 4'hD;
    SS2[18][44] = 4'hD;
    SS2[19][44] = 4'hC;
    SS2[20][44] = 4'hC;
    SS2[21][44] = 4'hC;
    SS2[22][44] = 4'hC;
    SS2[23][44] = 4'h0;
    SS2[24][44] = 4'h0;
    SS2[25][44] = 4'h0;
    SS2[26][44] = 4'h0;
    SS2[27][44] = 4'h0;
    SS2[28][44] = 4'h0;
    SS2[29][44] = 4'h0;
    SS2[30][44] = 4'h0;
    SS2[31][44] = 4'h0;
    SS2[32][44] = 4'hD;
    SS2[33][44] = 4'hD;
    SS2[34][44] = 4'hD;
    SS2[35][44] = 4'hD;
    SS2[36][44] = 4'h0;
    SS2[37][44] = 4'h0;
    SS2[38][44] = 4'h0;
    SS2[39][44] = 4'h0;
    SS2[40][44] = 4'h0;
    SS2[41][44] = 4'h0;
    SS2[42][44] = 4'h0;
    SS2[43][44] = 4'h0;
    SS2[44][44] = 4'h0;
    SS2[45][44] = 4'h0;
    SS2[46][44] = 4'h0;
    SS2[47][44] = 4'h0;
    SS2[0][45] = 4'h0;
    SS2[1][45] = 4'h0;
    SS2[2][45] = 4'h0;
    SS2[3][45] = 4'h0;
    SS2[4][45] = 4'h0;
    SS2[5][45] = 4'h0;
    SS2[6][45] = 4'h0;
    SS2[7][45] = 4'h0;
    SS2[8][45] = 4'h0;
    SS2[9][45] = 4'h0;
    SS2[10][45] = 4'h0;
    SS2[11][45] = 4'h0;
    SS2[12][45] = 4'h0;
    SS2[13][45] = 4'h0;
    SS2[14][45] = 4'h0;
    SS2[15][45] = 4'h0;
    SS2[16][45] = 4'hD;
    SS2[17][45] = 4'hD;
    SS2[18][45] = 4'hD;
    SS2[19][45] = 4'hC;
    SS2[20][45] = 4'hC;
    SS2[21][45] = 4'hC;
    SS2[22][45] = 4'hC;
    SS2[23][45] = 4'hC;
    SS2[24][45] = 4'h0;
    SS2[25][45] = 4'h0;
    SS2[26][45] = 4'h0;
    SS2[27][45] = 4'h0;
    SS2[28][45] = 4'h0;
    SS2[29][45] = 4'h0;
    SS2[30][45] = 4'h0;
    SS2[31][45] = 4'h0;
    SS2[32][45] = 4'h0;
    SS2[33][45] = 4'hD;
    SS2[34][45] = 4'hD;
    SS2[35][45] = 4'hD;
    SS2[36][45] = 4'h0;
    SS2[37][45] = 4'h0;
    SS2[38][45] = 4'h0;
    SS2[39][45] = 4'h0;
    SS2[40][45] = 4'h0;
    SS2[41][45] = 4'h0;
    SS2[42][45] = 4'h0;
    SS2[43][45] = 4'h0;
    SS2[44][45] = 4'h0;
    SS2[45][45] = 4'h0;
    SS2[46][45] = 4'h0;
    SS2[47][45] = 4'h0;
    SS2[0][46] = 4'h0;
    SS2[1][46] = 4'h0;
    SS2[2][46] = 4'h0;
    SS2[3][46] = 4'h0;
    SS2[4][46] = 4'h0;
    SS2[5][46] = 4'h0;
    SS2[6][46] = 4'h0;
    SS2[7][46] = 4'h0;
    SS2[8][46] = 4'h0;
    SS2[9][46] = 4'h0;
    SS2[10][46] = 4'h0;
    SS2[11][46] = 4'h0;
    SS2[12][46] = 4'h0;
    SS2[13][46] = 4'h0;
    SS2[14][46] = 4'h0;
    SS2[15][46] = 4'h0;
    SS2[16][46] = 4'h0;
    SS2[17][46] = 4'hD;
    SS2[18][46] = 4'hC;
    SS2[19][46] = 4'hC;
    SS2[20][46] = 4'hC;
    SS2[21][46] = 4'hC;
    SS2[22][46] = 4'hC;
    SS2[23][46] = 4'h0;
    SS2[24][46] = 4'h0;
    SS2[25][46] = 4'h0;
    SS2[26][46] = 4'h0;
    SS2[27][46] = 4'h0;
    SS2[28][46] = 4'h0;
    SS2[29][46] = 4'h0;
    SS2[30][46] = 4'h0;
    SS2[31][46] = 4'h0;
    SS2[32][46] = 4'h0;
    SS2[33][46] = 4'h0;
    SS2[34][46] = 4'hD;
    SS2[35][46] = 4'h0;
    SS2[36][46] = 4'h0;
    SS2[37][46] = 4'h0;
    SS2[38][46] = 4'h0;
    SS2[39][46] = 4'h0;
    SS2[40][46] = 4'h0;
    SS2[41][46] = 4'h0;
    SS2[42][46] = 4'h0;
    SS2[43][46] = 4'h0;
    SS2[44][46] = 4'h0;
    SS2[45][46] = 4'h0;
    SS2[46][46] = 4'h0;
    SS2[47][46] = 4'h0;
    SS2[0][47] = 4'h0;
    SS2[1][47] = 4'h0;
    SS2[2][47] = 4'h0;
    SS2[3][47] = 4'h0;
    SS2[4][47] = 4'h0;
    SS2[5][47] = 4'h0;
    SS2[6][47] = 4'h0;
    SS2[7][47] = 4'h0;
    SS2[8][47] = 4'h0;
    SS2[9][47] = 4'h0;
    SS2[10][47] = 4'h0;
    SS2[11][47] = 4'h0;
    SS2[12][47] = 4'h0;
    SS2[13][47] = 4'h0;
    SS2[14][47] = 4'h0;
    SS2[15][47] = 4'h0;
    SS2[16][47] = 4'h0;
    SS2[17][47] = 4'hE;
    SS2[18][47] = 4'hC;
    SS2[19][47] = 4'hC;
    SS2[20][47] = 4'hC;
    SS2[21][47] = 4'hC;
    SS2[22][47] = 4'h0;
    SS2[23][47] = 4'h0;
    SS2[24][47] = 4'h0;
    SS2[25][47] = 4'h0;
    SS2[26][47] = 4'h0;
    SS2[27][47] = 4'h0;
    SS2[28][47] = 4'h0;
    SS2[29][47] = 4'h0;
    SS2[30][47] = 4'h0;
    SS2[31][47] = 4'h0;
    SS2[32][47] = 4'h0;
    SS2[33][47] = 4'h0;
    SS2[34][47] = 4'h0;
    SS2[35][47] = 4'h0;
    SS2[36][47] = 4'h0;
    SS2[37][47] = 4'h0;
    SS2[38][47] = 4'h0;
    SS2[39][47] = 4'h0;
    SS2[40][47] = 4'h0;
    SS2[41][47] = 4'h0;
    SS2[42][47] = 4'h0;
    SS2[43][47] = 4'h0;
    SS2[44][47] = 4'h0;
    SS2[45][47] = 4'h0;
    SS2[46][47] = 4'h0;
    SS2[47][47] = 4'h0;
 
//SS 3
    SS3[0][0] = 4'h0;
    SS3[1][0] = 4'h0;
    SS3[2][0] = 4'h0;
    SS3[3][0] = 4'h0;
    SS3[4][0] = 4'h0;
    SS3[5][0] = 4'h0;
    SS3[6][0] = 4'h0;
    SS3[7][0] = 4'h0;
    SS3[8][0] = 4'h0;
    SS3[9][0] = 4'h0;
    SS3[10][0] = 4'h0;
    SS3[11][0] = 4'h0;
    SS3[12][0] = 4'h0;
    SS3[13][0] = 4'h0;
    SS3[14][0] = 4'h0;
    SS3[15][0] = 4'h0;
    SS3[16][0] = 4'h0;
    SS3[17][0] = 4'h0;
    SS3[18][0] = 4'h0;
    SS3[19][0] = 4'h0;
    SS3[20][0] = 4'h0;
    SS3[21][0] = 4'h0;
    SS3[22][0] = 4'h0;
    SS3[23][0] = 4'h0;
    SS3[24][0] = 4'h0;
    SS3[25][0] = 4'h0;
    SS3[26][0] = 4'h0;
    SS3[27][0] = 4'h0;
    SS3[28][0] = 4'h0;
    SS3[29][0] = 4'h0;
    SS3[30][0] = 4'h0;
    SS3[31][0] = 4'h0;
    SS3[32][0] = 4'h0;
    SS3[33][0] = 4'h0;
    SS3[34][0] = 4'h0;
    SS3[35][0] = 4'h0;
    SS3[36][0] = 4'h0;
    SS3[37][0] = 4'h0;
    SS3[38][0] = 4'h0;
    SS3[39][0] = 4'h0;
    SS3[40][0] = 4'h0;
    SS3[41][0] = 4'h0;
    SS3[42][0] = 4'h0;
    SS3[43][0] = 4'h0;
    SS3[44][0] = 4'h0;
    SS3[45][0] = 4'h0;
    SS3[46][0] = 4'h0;
    SS3[47][0] = 4'h0;
    SS3[0][1] = 4'h0;
    SS3[1][1] = 4'h0;
    SS3[2][1] = 4'h0;
    SS3[3][1] = 4'h0;
    SS3[4][1] = 4'h0;
    SS3[5][1] = 4'h0;
    SS3[6][1] = 4'h0;
    SS3[7][1] = 4'h0;
    SS3[8][1] = 4'h0;
    SS3[9][1] = 4'h0;
    SS3[10][1] = 4'h0;
    SS3[11][1] = 4'h0;
    SS3[12][1] = 4'h0;
    SS3[13][1] = 4'h0;
    SS3[14][1] = 4'h0;
    SS3[15][1] = 4'h0;
    SS3[16][1] = 4'h0;
    SS3[17][1] = 4'h0;
    SS3[18][1] = 4'h0;
    SS3[19][1] = 4'h0;
    SS3[20][1] = 4'h0;
    SS3[21][1] = 4'h0;
    SS3[22][1] = 4'h0;
    SS3[23][1] = 4'h0;
    SS3[24][1] = 4'h0;
    SS3[25][1] = 4'h0;
    SS3[26][1] = 4'h0;
    SS3[27][1] = 4'h0;
    SS3[28][1] = 4'h0;
    SS3[29][1] = 4'h0;
    SS3[30][1] = 4'h0;
    SS3[31][1] = 4'h0;
    SS3[32][1] = 4'h0;
    SS3[33][1] = 4'h0;
    SS3[34][1] = 4'h0;
    SS3[35][1] = 4'h0;
    SS3[36][1] = 4'h0;
    SS3[37][1] = 4'h0;
    SS3[38][1] = 4'h0;
    SS3[39][1] = 4'h0;
    SS3[40][1] = 4'h0;
    SS3[41][1] = 4'h0;
    SS3[42][1] = 4'h0;
    SS3[43][1] = 4'h0;
    SS3[44][1] = 4'h0;
    SS3[45][1] = 4'h0;
    SS3[46][1] = 4'h0;
    SS3[47][1] = 4'h0;
    SS3[0][2] = 4'h0;
    SS3[1][2] = 4'h0;
    SS3[2][2] = 4'h0;
    SS3[3][2] = 4'h0;
    SS3[4][2] = 4'h0;
    SS3[5][2] = 4'h0;
    SS3[6][2] = 4'h0;
    SS3[7][2] = 4'h0;
    SS3[8][2] = 4'h0;
    SS3[9][2] = 4'h0;
    SS3[10][2] = 4'h0;
    SS3[11][2] = 4'h0;
    SS3[12][2] = 4'h0;
    SS3[13][2] = 4'h0;
    SS3[14][2] = 4'h0;
    SS3[15][2] = 4'h0;
    SS3[16][2] = 4'h0;
    SS3[17][2] = 4'h0;
    SS3[18][2] = 4'h0;
    SS3[19][2] = 4'h0;
    SS3[20][2] = 4'h0;
    SS3[21][2] = 4'h0;
    SS3[22][2] = 4'h0;
    SS3[23][2] = 4'h0;
    SS3[24][2] = 4'h0;
    SS3[25][2] = 4'h0;
    SS3[26][2] = 4'h0;
    SS3[27][2] = 4'h0;
    SS3[28][2] = 4'h0;
    SS3[29][2] = 4'h0;
    SS3[30][2] = 4'h0;
    SS3[31][2] = 4'h0;
    SS3[32][2] = 4'h0;
    SS3[33][2] = 4'h0;
    SS3[34][2] = 4'h0;
    SS3[35][2] = 4'h0;
    SS3[36][2] = 4'h0;
    SS3[37][2] = 4'h0;
    SS3[38][2] = 4'h0;
    SS3[39][2] = 4'h0;
    SS3[40][2] = 4'h0;
    SS3[41][2] = 4'h0;
    SS3[42][2] = 4'h0;
    SS3[43][2] = 4'h0;
    SS3[44][2] = 4'h0;
    SS3[45][2] = 4'h0;
    SS3[46][2] = 4'h0;
    SS3[47][2] = 4'h0;
    SS3[0][3] = 4'h0;
    SS3[1][3] = 4'h0;
    SS3[2][3] = 4'h0;
    SS3[3][3] = 4'h0;
    SS3[4][3] = 4'h0;
    SS3[5][3] = 4'h0;
    SS3[6][3] = 4'h0;
    SS3[7][3] = 4'h0;
    SS3[8][3] = 4'h0;
    SS3[9][3] = 4'h0;
    SS3[10][3] = 4'h0;
    SS3[11][3] = 4'h0;
    SS3[12][3] = 4'h0;
    SS3[13][3] = 4'h0;
    SS3[14][3] = 4'h0;
    SS3[15][3] = 4'h0;
    SS3[16][3] = 4'h0;
    SS3[17][3] = 4'h0;
    SS3[18][3] = 4'h0;
    SS3[19][3] = 4'h0;
    SS3[20][3] = 4'h0;
    SS3[21][3] = 4'h0;
    SS3[22][3] = 4'h0;
    SS3[23][3] = 4'h0;
    SS3[24][3] = 4'h0;
    SS3[25][3] = 4'h0;
    SS3[26][3] = 4'h0;
    SS3[27][3] = 4'h0;
    SS3[28][3] = 4'h0;
    SS3[29][3] = 4'h0;
    SS3[30][3] = 4'h0;
    SS3[31][3] = 4'h0;
    SS3[32][3] = 4'h0;
    SS3[33][3] = 4'h0;
    SS3[34][3] = 4'h0;
    SS3[35][3] = 4'h0;
    SS3[36][3] = 4'h0;
    SS3[37][3] = 4'h0;
    SS3[38][3] = 4'h0;
    SS3[39][3] = 4'h0;
    SS3[40][3] = 4'h0;
    SS3[41][3] = 4'h0;
    SS3[42][3] = 4'h0;
    SS3[43][3] = 4'h0;
    SS3[44][3] = 4'h0;
    SS3[45][3] = 4'h0;
    SS3[46][3] = 4'h0;
    SS3[47][3] = 4'h0;
    SS3[0][4] = 4'h0;
    SS3[1][4] = 4'h0;
    SS3[2][4] = 4'h0;
    SS3[3][4] = 4'h0;
    SS3[4][4] = 4'h0;
    SS3[5][4] = 4'h0;
    SS3[6][4] = 4'h0;
    SS3[7][4] = 4'h0;
    SS3[8][4] = 4'h0;
    SS3[9][4] = 4'hD;
    SS3[10][4] = 4'h0;
    SS3[11][4] = 4'h0;
    SS3[12][4] = 4'h0;
    SS3[13][4] = 4'h0;
    SS3[14][4] = 4'h0;
    SS3[15][4] = 4'h0;
    SS3[16][4] = 4'h0;
    SS3[17][4] = 4'h0;
    SS3[18][4] = 4'h0;
    SS3[19][4] = 4'h0;
    SS3[20][4] = 4'h0;
    SS3[21][4] = 4'h0;
    SS3[22][4] = 4'h0;
    SS3[23][4] = 4'h0;
    SS3[24][4] = 4'h0;
    SS3[25][4] = 4'h0;
    SS3[26][4] = 4'h0;
    SS3[27][4] = 4'h0;
    SS3[28][4] = 4'h0;
    SS3[29][4] = 4'h0;
    SS3[30][4] = 4'h0;
    SS3[31][4] = 4'h0;
    SS3[32][4] = 4'h0;
    SS3[33][4] = 4'h0;
    SS3[34][4] = 4'h0;
    SS3[35][4] = 4'h0;
    SS3[36][4] = 4'h0;
    SS3[37][4] = 4'h0;
    SS3[38][4] = 4'h0;
    SS3[39][4] = 4'h0;
    SS3[40][4] = 4'h0;
    SS3[41][4] = 4'h0;
    SS3[42][4] = 4'h0;
    SS3[43][4] = 4'h0;
    SS3[44][4] = 4'h0;
    SS3[45][4] = 4'h0;
    SS3[46][4] = 4'h0;
    SS3[47][4] = 4'h0;
    SS3[0][5] = 4'h0;
    SS3[1][5] = 4'h0;
    SS3[2][5] = 4'h0;
    SS3[3][5] = 4'h0;
    SS3[4][5] = 4'h0;
    SS3[5][5] = 4'h0;
    SS3[6][5] = 4'h0;
    SS3[7][5] = 4'hD;
    SS3[8][5] = 4'hD;
    SS3[9][5] = 4'hD;
    SS3[10][5] = 4'h0;
    SS3[11][5] = 4'h0;
    SS3[12][5] = 4'h0;
    SS3[13][5] = 4'h0;
    SS3[14][5] = 4'h0;
    SS3[15][5] = 4'h0;
    SS3[16][5] = 4'h0;
    SS3[17][5] = 4'h0;
    SS3[18][5] = 4'h0;
    SS3[19][5] = 4'h0;
    SS3[20][5] = 4'h0;
    SS3[21][5] = 4'h0;
    SS3[22][5] = 4'h0;
    SS3[23][5] = 4'h0;
    SS3[24][5] = 4'h0;
    SS3[25][5] = 4'h0;
    SS3[26][5] = 4'h0;
    SS3[27][5] = 4'h0;
    SS3[28][5] = 4'h0;
    SS3[29][5] = 4'h0;
    SS3[30][5] = 4'h0;
    SS3[31][5] = 4'h0;
    SS3[32][5] = 4'h0;
    SS3[33][5] = 4'h0;
    SS3[34][5] = 4'h0;
    SS3[35][5] = 4'h0;
    SS3[36][5] = 4'h0;
    SS3[37][5] = 4'h0;
    SS3[38][5] = 4'h0;
    SS3[39][5] = 4'h0;
    SS3[40][5] = 4'h0;
    SS3[41][5] = 4'h0;
    SS3[42][5] = 4'h0;
    SS3[43][5] = 4'h0;
    SS3[44][5] = 4'h0;
    SS3[45][5] = 4'h0;
    SS3[46][5] = 4'h0;
    SS3[47][5] = 4'h0;
    SS3[0][6] = 4'h0;
    SS3[1][6] = 4'h0;
    SS3[2][6] = 4'h0;
    SS3[3][6] = 4'h0;
    SS3[4][6] = 4'h0;
    SS3[5][6] = 4'h0;
    SS3[6][6] = 4'h0;
    SS3[7][6] = 4'hD;
    SS3[8][6] = 4'hD;
    SS3[9][6] = 4'hD;
    SS3[10][6] = 4'h0;
    SS3[11][6] = 4'h0;
    SS3[12][6] = 4'hD;
    SS3[13][6] = 4'hD;
    SS3[14][6] = 4'h0;
    SS3[15][6] = 4'h0;
    SS3[16][6] = 4'h0;
    SS3[17][6] = 4'h0;
    SS3[18][6] = 4'h0;
    SS3[19][6] = 4'h0;
    SS3[20][6] = 4'h0;
    SS3[21][6] = 4'h0;
    SS3[22][6] = 4'h0;
    SS3[23][6] = 4'h0;
    SS3[24][6] = 4'h0;
    SS3[25][6] = 4'h0;
    SS3[26][6] = 4'h0;
    SS3[27][6] = 4'h0;
    SS3[28][6] = 4'h0;
    SS3[29][6] = 4'h0;
    SS3[30][6] = 4'h0;
    SS3[31][6] = 4'h0;
    SS3[32][6] = 4'h0;
    SS3[33][6] = 4'h0;
    SS3[34][6] = 4'h0;
    SS3[35][6] = 4'h0;
    SS3[36][6] = 4'h0;
    SS3[37][6] = 4'h0;
    SS3[38][6] = 4'h0;
    SS3[39][6] = 4'h0;
    SS3[40][6] = 4'h0;
    SS3[41][6] = 4'h0;
    SS3[42][6] = 4'h0;
    SS3[43][6] = 4'h0;
    SS3[44][6] = 4'h0;
    SS3[45][6] = 4'h0;
    SS3[46][6] = 4'h0;
    SS3[47][6] = 4'h0;
    SS3[0][7] = 4'h0;
    SS3[1][7] = 4'h0;
    SS3[2][7] = 4'h0;
    SS3[3][7] = 4'h0;
    SS3[4][7] = 4'h0;
    SS3[5][7] = 4'h0;
    SS3[6][7] = 4'h0;
    SS3[7][7] = 4'h0;
    SS3[8][7] = 4'hD;
    SS3[9][7] = 4'hD;
    SS3[10][7] = 4'hD;
    SS3[11][7] = 4'hD;
    SS3[12][7] = 4'hD;
    SS3[13][7] = 4'hD;
    SS3[14][7] = 4'h0;
    SS3[15][7] = 4'h0;
    SS3[16][7] = 4'h0;
    SS3[17][7] = 4'h0;
    SS3[18][7] = 4'h0;
    SS3[19][7] = 4'h0;
    SS3[20][7] = 4'h0;
    SS3[21][7] = 4'h0;
    SS3[22][7] = 4'h0;
    SS3[23][7] = 4'h0;
    SS3[24][7] = 4'h0;
    SS3[25][7] = 4'h0;
    SS3[26][7] = 4'h0;
    SS3[27][7] = 4'h0;
    SS3[28][7] = 4'h0;
    SS3[29][7] = 4'h0;
    SS3[30][7] = 4'h0;
    SS3[31][7] = 4'h0;
    SS3[32][7] = 4'h0;
    SS3[33][7] = 4'h0;
    SS3[34][7] = 4'h0;
    SS3[35][7] = 4'h0;
    SS3[36][7] = 4'h0;
    SS3[37][7] = 4'h0;
    SS3[38][7] = 4'h0;
    SS3[39][7] = 4'h0;
    SS3[40][7] = 4'h0;
    SS3[41][7] = 4'h0;
    SS3[42][7] = 4'h0;
    SS3[43][7] = 4'h0;
    SS3[44][7] = 4'h0;
    SS3[45][7] = 4'h0;
    SS3[46][7] = 4'h0;
    SS3[47][7] = 4'h0;
    SS3[0][8] = 4'h0;
    SS3[1][8] = 4'h0;
    SS3[2][8] = 4'h0;
    SS3[3][8] = 4'h0;
    SS3[4][8] = 4'h0;
    SS3[5][8] = 4'h0;
    SS3[6][8] = 4'h0;
    SS3[7][8] = 4'h0;
    SS3[8][8] = 4'hD;
    SS3[9][8] = 4'hD;
    SS3[10][8] = 4'hD;
    SS3[11][8] = 4'hD;
    SS3[12][8] = 4'hD;
    SS3[13][8] = 4'hD;
    SS3[14][8] = 4'h0;
    SS3[15][8] = 4'h3;
    SS3[16][8] = 4'h3;
    SS3[17][8] = 4'h3;
    SS3[18][8] = 4'h0;
    SS3[19][8] = 4'h0;
    SS3[20][8] = 4'h0;
    SS3[21][8] = 4'h0;
    SS3[22][8] = 4'h0;
    SS3[23][8] = 4'h0;
    SS3[24][8] = 4'h0;
    SS3[25][8] = 4'h0;
    SS3[26][8] = 4'h0;
    SS3[27][8] = 4'h0;
    SS3[28][8] = 4'h0;
    SS3[29][8] = 4'h0;
    SS3[30][8] = 4'h0;
    SS3[31][8] = 4'h0;
    SS3[32][8] = 4'h0;
    SS3[33][8] = 4'h0;
    SS3[34][8] = 4'h0;
    SS3[35][8] = 4'h0;
    SS3[36][8] = 4'h0;
    SS3[37][8] = 4'h0;
    SS3[38][8] = 4'h0;
    SS3[39][8] = 4'h0;
    SS3[40][8] = 4'h0;
    SS3[41][8] = 4'h0;
    SS3[42][8] = 4'h0;
    SS3[43][8] = 4'h0;
    SS3[44][8] = 4'h0;
    SS3[45][8] = 4'h0;
    SS3[46][8] = 4'h0;
    SS3[47][8] = 4'h0;
    SS3[0][9] = 4'h0;
    SS3[1][9] = 4'h0;
    SS3[2][9] = 4'h0;
    SS3[3][9] = 4'h0;
    SS3[4][9] = 4'h0;
    SS3[5][9] = 4'h0;
    SS3[6][9] = 4'h0;
    SS3[7][9] = 4'h0;
    SS3[8][9] = 4'hD;
    SS3[9][9] = 4'hD;
    SS3[10][9] = 4'hD;
    SS3[11][9] = 4'hD;
    SS3[12][9] = 4'hD;
    SS3[13][9] = 4'hD;
    SS3[14][9] = 4'hD;
    SS3[15][9] = 4'h3;
    SS3[16][9] = 4'h3;
    SS3[17][9] = 4'h3;
    SS3[18][9] = 4'h0;
    SS3[19][9] = 4'h0;
    SS3[20][9] = 4'h0;
    SS3[21][9] = 4'h0;
    SS3[22][9] = 4'h0;
    SS3[23][9] = 4'h0;
    SS3[24][9] = 4'h0;
    SS3[25][9] = 4'h0;
    SS3[26][9] = 4'h0;
    SS3[27][9] = 4'h0;
    SS3[28][9] = 4'h0;
    SS3[29][9] = 4'h0;
    SS3[30][9] = 4'h0;
    SS3[31][9] = 4'h0;
    SS3[32][9] = 4'h0;
    SS3[33][9] = 4'h0;
    SS3[34][9] = 4'h0;
    SS3[35][9] = 4'h0;
    SS3[36][9] = 4'h0;
    SS3[37][9] = 4'h0;
    SS3[38][9] = 4'h0;
    SS3[39][9] = 4'h0;
    SS3[40][9] = 4'h0;
    SS3[41][9] = 4'h0;
    SS3[42][9] = 4'h0;
    SS3[43][9] = 4'h0;
    SS3[44][9] = 4'h0;
    SS3[45][9] = 4'h0;
    SS3[46][9] = 4'h0;
    SS3[47][9] = 4'h0;
    SS3[0][10] = 4'h0;
    SS3[1][10] = 4'h0;
    SS3[2][10] = 4'h0;
    SS3[3][10] = 4'h0;
    SS3[4][10] = 4'h0;
    SS3[5][10] = 4'h0;
    SS3[6][10] = 4'h0;
    SS3[7][10] = 4'h0;
    SS3[8][10] = 4'h0;
    SS3[9][10] = 4'hD;
    SS3[10][10] = 4'hE;
    SS3[11][10] = 4'hE;
    SS3[12][10] = 4'hD;
    SS3[13][10] = 4'hD;
    SS3[14][10] = 4'hD;
    SS3[15][10] = 4'h3;
    SS3[16][10] = 4'h3;
    SS3[17][10] = 4'h3;
    SS3[18][10] = 4'h0;
    SS3[19][10] = 4'h0;
    SS3[20][10] = 4'h0;
    SS3[21][10] = 4'h0;
    SS3[22][10] = 4'h0;
    SS3[23][10] = 4'h0;
    SS3[24][10] = 4'h0;
    SS3[25][10] = 4'h0;
    SS3[26][10] = 4'h0;
    SS3[27][10] = 4'h0;
    SS3[28][10] = 4'h0;
    SS3[29][10] = 4'h0;
    SS3[30][10] = 4'h0;
    SS3[31][10] = 4'h0;
    SS3[32][10] = 4'h0;
    SS3[33][10] = 4'h0;
    SS3[34][10] = 4'h0;
    SS3[35][10] = 4'h0;
    SS3[36][10] = 4'h0;
    SS3[37][10] = 4'h0;
    SS3[38][10] = 4'h0;
    SS3[39][10] = 4'h0;
    SS3[40][10] = 4'h0;
    SS3[41][10] = 4'h0;
    SS3[42][10] = 4'h0;
    SS3[43][10] = 4'h0;
    SS3[44][10] = 4'h0;
    SS3[45][10] = 4'h0;
    SS3[46][10] = 4'h0;
    SS3[47][10] = 4'h0;
    SS3[0][11] = 4'h0;
    SS3[1][11] = 4'h0;
    SS3[2][11] = 4'h0;
    SS3[3][11] = 4'h0;
    SS3[4][11] = 4'h0;
    SS3[5][11] = 4'h0;
    SS3[6][11] = 4'h0;
    SS3[7][11] = 4'h0;
    SS3[8][11] = 4'h0;
    SS3[9][11] = 4'hE;
    SS3[10][11] = 4'hE;
    SS3[11][11] = 4'hE;
    SS3[12][11] = 4'hD;
    SS3[13][11] = 4'hD;
    SS3[14][11] = 4'hD;
    SS3[15][11] = 4'hE;
    SS3[16][11] = 4'hD;
    SS3[17][11] = 4'hD;
    SS3[18][11] = 4'hD;
    SS3[19][11] = 4'h0;
    SS3[20][11] = 4'h0;
    SS3[21][11] = 4'h0;
    SS3[22][11] = 4'h0;
    SS3[23][11] = 4'h3;
    SS3[24][11] = 4'h3;
    SS3[25][11] = 4'h0;
    SS3[26][11] = 4'h0;
    SS3[27][11] = 4'h0;
    SS3[28][11] = 4'h0;
    SS3[29][11] = 4'h0;
    SS3[30][11] = 4'h0;
    SS3[31][11] = 4'h0;
    SS3[32][11] = 4'h0;
    SS3[33][11] = 4'h0;
    SS3[34][11] = 4'h0;
    SS3[35][11] = 4'h0;
    SS3[36][11] = 4'h0;
    SS3[37][11] = 4'h0;
    SS3[38][11] = 4'h0;
    SS3[39][11] = 4'h0;
    SS3[40][11] = 4'h0;
    SS3[41][11] = 4'h0;
    SS3[42][11] = 4'h0;
    SS3[43][11] = 4'h0;
    SS3[44][11] = 4'h0;
    SS3[45][11] = 4'h0;
    SS3[46][11] = 4'h0;
    SS3[47][11] = 4'h0;
    SS3[0][12] = 4'h0;
    SS3[1][12] = 4'h0;
    SS3[2][12] = 4'h0;
    SS3[3][12] = 4'h0;
    SS3[4][12] = 4'h0;
    SS3[5][12] = 4'h0;
    SS3[6][12] = 4'h0;
    SS3[7][12] = 4'h0;
    SS3[8][12] = 4'h0;
    SS3[9][12] = 4'h0;
    SS3[10][12] = 4'hE;
    SS3[11][12] = 4'hE;
    SS3[12][12] = 4'hE;
    SS3[13][12] = 4'hE;
    SS3[14][12] = 4'hE;
    SS3[15][12] = 4'hE;
    SS3[16][12] = 4'hD;
    SS3[17][12] = 4'hD;
    SS3[18][12] = 4'hD;
    SS3[19][12] = 4'h0;
    SS3[20][12] = 4'h0;
    SS3[21][12] = 4'hD;
    SS3[22][12] = 4'h3;
    SS3[23][12] = 4'h3;
    SS3[24][12] = 4'h3;
    SS3[25][12] = 4'h3;
    SS3[26][12] = 4'h0;
    SS3[27][12] = 4'h0;
    SS3[28][12] = 4'h0;
    SS3[29][12] = 4'h0;
    SS3[30][12] = 4'h0;
    SS3[31][12] = 4'h0;
    SS3[32][12] = 4'h0;
    SS3[33][12] = 4'h0;
    SS3[34][12] = 4'h0;
    SS3[35][12] = 4'h0;
    SS3[36][12] = 4'hD;
    SS3[37][12] = 4'hD;
    SS3[38][12] = 4'hF;
    SS3[39][12] = 4'h0;
    SS3[40][12] = 4'h0;
    SS3[41][12] = 4'h0;
    SS3[42][12] = 4'h0;
    SS3[43][12] = 4'h0;
    SS3[44][12] = 4'hC;
    SS3[45][12] = 4'h0;
    SS3[46][12] = 4'h0;
    SS3[47][12] = 4'h0;
    SS3[0][13] = 4'h0;
    SS3[1][13] = 4'h0;
    SS3[2][13] = 4'h0;
    SS3[3][13] = 4'h0;
    SS3[4][13] = 4'h0;
    SS3[5][13] = 4'h0;
    SS3[6][13] = 4'h0;
    SS3[7][13] = 4'h0;
    SS3[8][13] = 4'h0;
    SS3[9][13] = 4'h0;
    SS3[10][13] = 4'hE;
    SS3[11][13] = 4'hE;
    SS3[12][13] = 4'hE;
    SS3[13][13] = 4'hE;
    SS3[14][13] = 4'hE;
    SS3[15][13] = 4'hE;
    SS3[16][13] = 4'hD;
    SS3[17][13] = 4'hD;
    SS3[18][13] = 4'hD;
    SS3[19][13] = 4'hD;
    SS3[20][13] = 4'hD;
    SS3[21][13] = 4'hD;
    SS3[22][13] = 4'hD;
    SS3[23][13] = 4'h3;
    SS3[24][13] = 4'h3;
    SS3[25][13] = 4'h3;
    SS3[26][13] = 4'h0;
    SS3[27][13] = 4'h0;
    SS3[28][13] = 4'h0;
    SS3[29][13] = 4'h0;
    SS3[30][13] = 4'h0;
    SS3[31][13] = 4'h0;
    SS3[32][13] = 4'h0;
    SS3[33][13] = 4'h0;
    SS3[34][13] = 4'hD;
    SS3[35][13] = 4'hD;
    SS3[36][13] = 4'hD;
    SS3[37][13] = 4'hD;
    SS3[38][13] = 4'hD;
    SS3[39][13] = 4'h0;
    SS3[40][13] = 4'h0;
    SS3[41][13] = 4'h0;
    SS3[42][13] = 4'hC;
    SS3[43][13] = 4'hC;
    SS3[44][13] = 4'hC;
    SS3[45][13] = 4'h0;
    SS3[46][13] = 4'h0;
    SS3[47][13] = 4'h0;
    SS3[0][14] = 4'h0;
    SS3[1][14] = 4'h0;
    SS3[2][14] = 4'h0;
    SS3[3][14] = 4'h0;
    SS3[4][14] = 4'h0;
    SS3[5][14] = 4'h0;
    SS3[6][14] = 4'h0;
    SS3[7][14] = 4'h0;
    SS3[8][14] = 4'h0;
    SS3[9][14] = 4'h0;
    SS3[10][14] = 4'hE;
    SS3[11][14] = 4'hE;
    SS3[12][14] = 4'hE;
    SS3[13][14] = 4'hE;
    SS3[14][14] = 4'hE;
    SS3[15][14] = 4'hE;
    SS3[16][14] = 4'hE;
    SS3[17][14] = 4'hD;
    SS3[18][14] = 4'hD;
    SS3[19][14] = 4'hD;
    SS3[20][14] = 4'hD;
    SS3[21][14] = 4'hD;
    SS3[22][14] = 4'hD;
    SS3[23][14] = 4'h3;
    SS3[24][14] = 4'hD;
    SS3[25][14] = 4'hD;
    SS3[26][14] = 4'hF;
    SS3[27][14] = 4'h0;
    SS3[28][14] = 4'h0;
    SS3[29][14] = 4'h0;
    SS3[30][14] = 4'h0;
    SS3[31][14] = 4'hD;
    SS3[32][14] = 4'hD;
    SS3[33][14] = 4'hD;
    SS3[34][14] = 4'hD;
    SS3[35][14] = 4'hD;
    SS3[36][14] = 4'hD;
    SS3[37][14] = 4'hD;
    SS3[38][14] = 4'hD;
    SS3[39][14] = 4'hC;
    SS3[40][14] = 4'hC;
    SS3[41][14] = 4'hC;
    SS3[42][14] = 4'hC;
    SS3[43][14] = 4'hC;
    SS3[44][14] = 4'hC;
    SS3[45][14] = 4'hC;
    SS3[46][14] = 4'h0;
    SS3[47][14] = 4'h0;
    SS3[0][15] = 4'h0;
    SS3[1][15] = 4'h0;
    SS3[2][15] = 4'h0;
    SS3[3][15] = 4'h0;
    SS3[4][15] = 4'h0;
    SS3[5][15] = 4'h0;
    SS3[6][15] = 4'h0;
    SS3[7][15] = 4'h0;
    SS3[8][15] = 4'h0;
    SS3[9][15] = 4'h0;
    SS3[10][15] = 4'h0;
    SS3[11][15] = 4'hE;
    SS3[12][15] = 4'hE;
    SS3[13][15] = 4'hE;
    SS3[14][15] = 4'hE;
    SS3[15][15] = 4'hE;
    SS3[16][15] = 4'hE;
    SS3[17][15] = 4'hD;
    SS3[18][15] = 4'hD;
    SS3[19][15] = 4'hD;
    SS3[20][15] = 4'hD;
    SS3[21][15] = 4'hD;
    SS3[22][15] = 4'hD;
    SS3[23][15] = 4'hD;
    SS3[24][15] = 4'hD;
    SS3[25][15] = 4'hD;
    SS3[26][15] = 4'hD;
    SS3[27][15] = 4'h0;
    SS3[28][15] = 4'h0;
    SS3[29][15] = 4'hC;
    SS3[30][15] = 4'hD;
    SS3[31][15] = 4'hD;
    SS3[32][15] = 4'hD;
    SS3[33][15] = 4'hD;
    SS3[34][15] = 4'hD;
    SS3[35][15] = 4'hD;
    SS3[36][15] = 4'hD;
    SS3[37][15] = 4'hC;
    SS3[38][15] = 4'hC;
    SS3[39][15] = 4'hC;
    SS3[40][15] = 4'hC;
    SS3[41][15] = 4'hC;
    SS3[42][15] = 4'hC;
    SS3[43][15] = 4'hC;
    SS3[44][15] = 4'hC;
    SS3[45][15] = 4'hC;
    SS3[46][15] = 4'h0;
    SS3[47][15] = 4'h0;
    SS3[0][16] = 4'h0;
    SS3[1][16] = 4'h0;
    SS3[2][16] = 4'h0;
    SS3[3][16] = 4'hC;
    SS3[4][16] = 4'hC;
    SS3[5][16] = 4'h0;
    SS3[6][16] = 4'h0;
    SS3[7][16] = 4'h0;
    SS3[8][16] = 4'h0;
    SS3[9][16] = 4'h0;
    SS3[10][16] = 4'h0;
    SS3[11][16] = 4'hC;
    SS3[12][16] = 4'hC;
    SS3[13][16] = 4'hC;
    SS3[14][16] = 4'hE;
    SS3[15][16] = 4'hE;
    SS3[16][16] = 4'hE;
    SS3[17][16] = 4'hE;
    SS3[18][16] = 4'hD;
    SS3[19][16] = 4'hE;
    SS3[20][16] = 4'hE;
    SS3[21][16] = 4'hD;
    SS3[22][16] = 4'hD;
    SS3[23][16] = 4'hD;
    SS3[24][16] = 4'hD;
    SS3[25][16] = 4'hD;
    SS3[26][16] = 4'hD;
    SS3[27][16] = 4'hC;
    SS3[28][16] = 4'hC;
    SS3[29][16] = 4'hC;
    SS3[30][16] = 4'hC;
    SS3[31][16] = 4'hD;
    SS3[32][16] = 4'hD;
    SS3[33][16] = 4'hD;
    SS3[34][16] = 4'hC;
    SS3[35][16] = 4'hC;
    SS3[36][16] = 4'hC;
    SS3[37][16] = 4'hC;
    SS3[38][16] = 4'hC;
    SS3[39][16] = 4'hC;
    SS3[40][16] = 4'hC;
    SS3[41][16] = 4'hC;
    SS3[42][16] = 4'hC;
    SS3[43][16] = 4'hC;
    SS3[44][16] = 4'hC;
    SS3[45][16] = 4'hC;
    SS3[46][16] = 4'hC;
    SS3[47][16] = 4'h0;
    SS3[0][17] = 4'h0;
    SS3[1][17] = 4'hC;
    SS3[2][17] = 4'hC;
    SS3[3][17] = 4'hC;
    SS3[4][17] = 4'hC;
    SS3[5][17] = 4'h0;
    SS3[6][17] = 4'h0;
    SS3[7][17] = 4'h0;
    SS3[8][17] = 4'h0;
    SS3[9][17] = 4'hC;
    SS3[10][17] = 4'hC;
    SS3[11][17] = 4'hC;
    SS3[12][17] = 4'hC;
    SS3[13][17] = 4'hC;
    SS3[14][17] = 4'hC;
    SS3[15][17] = 4'hE;
    SS3[16][17] = 4'hC;
    SS3[17][17] = 4'hC;
    SS3[18][17] = 4'hE;
    SS3[19][17] = 4'hE;
    SS3[20][17] = 4'hE;
    SS3[21][17] = 4'hD;
    SS3[22][17] = 4'hD;
    SS3[23][17] = 4'hD;
    SS3[24][17] = 4'hC;
    SS3[25][17] = 4'hD;
    SS3[26][17] = 4'hD;
    SS3[27][17] = 4'hD;
    SS3[28][17] = 4'hC;
    SS3[29][17] = 4'hC;
    SS3[30][17] = 4'hC;
    SS3[31][17] = 4'hD;
    SS3[32][17] = 4'hC;
    SS3[33][17] = 4'hC;
    SS3[34][17] = 4'hC;
    SS3[35][17] = 4'hC;
    SS3[36][17] = 4'hC;
    SS3[37][17] = 4'hC;
    SS3[38][17] = 4'hC;
    SS3[39][17] = 4'hC;
    SS3[40][17] = 4'hC;
    SS3[41][17] = 4'hC;
    SS3[42][17] = 4'hC;
    SS3[43][17] = 4'hC;
    SS3[44][17] = 4'hC;
    SS3[45][17] = 4'hC;
    SS3[46][17] = 4'hC;
    SS3[47][17] = 4'h0;
    SS3[0][18] = 4'hC;
    SS3[1][18] = 4'hC;
    SS3[2][18] = 4'hC;
    SS3[3][18] = 4'hC;
    SS3[4][18] = 4'hC;
    SS3[5][18] = 4'hC;
    SS3[6][18] = 4'hC;
    SS3[7][18] = 4'hC;
    SS3[8][18] = 4'hC;
    SS3[9][18] = 4'hC;
    SS3[10][18] = 4'hC;
    SS3[11][18] = 4'hC;
    SS3[12][18] = 4'hC;
    SS3[13][18] = 4'hC;
    SS3[14][18] = 4'hC;
    SS3[15][18] = 4'hC;
    SS3[16][18] = 4'hC;
    SS3[17][18] = 4'hC;
    SS3[18][18] = 4'hC;
    SS3[19][18] = 4'hE;
    SS3[20][18] = 4'hE;
    SS3[21][18] = 4'hE;
    SS3[22][18] = 4'hC;
    SS3[23][18] = 4'hC;
    SS3[24][18] = 4'hC;
    SS3[25][18] = 4'hD;
    SS3[26][18] = 4'hD;
    SS3[27][18] = 4'hD;
    SS3[28][18] = 4'hC;
    SS3[29][18] = 4'hC;
    SS3[30][18] = 4'hC;
    SS3[31][18] = 4'hC;
    SS3[32][18] = 4'hC;
    SS3[33][18] = 4'hC;
    SS3[34][18] = 4'hC;
    SS3[35][18] = 4'hC;
    SS3[36][18] = 4'hC;
    SS3[37][18] = 4'hC;
    SS3[38][18] = 4'hC;
    SS3[39][18] = 4'hC;
    SS3[40][18] = 4'hC;
    SS3[41][18] = 4'hC;
    SS3[42][18] = 4'hC;
    SS3[43][18] = 4'hC;
    SS3[44][18] = 4'hC;
    SS3[45][18] = 4'h0;
    SS3[46][18] = 4'h0;
    SS3[47][18] = 4'h0;
    SS3[0][19] = 4'hC;
    SS3[1][19] = 4'hC;
    SS3[2][19] = 4'hC;
    SS3[3][19] = 4'hC;
    SS3[4][19] = 4'hC;
    SS3[5][19] = 4'hC;
    SS3[6][19] = 4'hC;
    SS3[7][19] = 4'hC;
    SS3[8][19] = 4'hC;
    SS3[9][19] = 4'hC;
    SS3[10][19] = 4'hC;
    SS3[11][19] = 4'hC;
    SS3[12][19] = 4'hC;
    SS3[13][19] = 4'hC;
    SS3[14][19] = 4'hC;
    SS3[15][19] = 4'hC;
    SS3[16][19] = 4'hC;
    SS3[17][19] = 4'hC;
    SS3[18][19] = 4'hC;
    SS3[19][19] = 4'hC;
    SS3[20][19] = 4'hC;
    SS3[21][19] = 4'hC;
    SS3[22][19] = 4'hC;
    SS3[23][19] = 4'hC;
    SS3[24][19] = 4'hC;
    SS3[25][19] = 4'hD;
    SS3[26][19] = 4'hD;
    SS3[27][19] = 4'hA;
    SS3[28][19] = 4'hA;
    SS3[29][19] = 4'hC;
    SS3[30][19] = 4'hC;
    SS3[31][19] = 4'hC;
    SS3[32][19] = 4'hC;
    SS3[33][19] = 4'hC;
    SS3[34][19] = 4'hC;
    SS3[35][19] = 4'hC;
    SS3[36][19] = 4'hC;
    SS3[37][19] = 4'hC;
    SS3[38][19] = 4'hC;
    SS3[39][19] = 4'hC;
    SS3[40][19] = 4'hC;
    SS3[41][19] = 4'hC;
    SS3[42][19] = 4'hC;
    SS3[43][19] = 4'h0;
    SS3[44][19] = 4'h0;
    SS3[45][19] = 4'h0;
    SS3[46][19] = 4'h0;
    SS3[47][19] = 4'h0;
    SS3[0][20] = 4'hC;
    SS3[1][20] = 4'hD;
    SS3[2][20] = 4'hD;
    SS3[3][20] = 4'hC;
    SS3[4][20] = 4'hC;
    SS3[5][20] = 4'hC;
    SS3[6][20] = 4'hC;
    SS3[7][20] = 4'hC;
    SS3[8][20] = 4'hC;
    SS3[9][20] = 4'hD;
    SS3[10][20] = 4'hC;
    SS3[11][20] = 4'hC;
    SS3[12][20] = 4'hC;
    SS3[13][20] = 4'hC;
    SS3[14][20] = 4'hC;
    SS3[15][20] = 4'hC;
    SS3[16][20] = 4'hC;
    SS3[17][20] = 4'hC;
    SS3[18][20] = 4'hC;
    SS3[19][20] = 4'hC;
    SS3[20][20] = 4'hC;
    SS3[21][20] = 4'hC;
    SS3[22][20] = 4'hC;
    SS3[23][20] = 4'hC;
    SS3[24][20] = 4'hC;
    SS3[25][20] = 4'hD;
    SS3[26][20] = 4'hA;
    SS3[27][20] = 4'hA;
    SS3[28][20] = 4'hA;
    SS3[29][20] = 4'hC;
    SS3[30][20] = 4'hC;
    SS3[31][20] = 4'hC;
    SS3[32][20] = 4'hC;
    SS3[33][20] = 4'hC;
    SS3[34][20] = 4'hC;
    SS3[35][20] = 4'hC;
    SS3[36][20] = 4'hC;
    SS3[37][20] = 4'hC;
    SS3[38][20] = 4'hC;
    SS3[39][20] = 4'hC;
    SS3[40][20] = 4'hD;
    SS3[41][20] = 4'hD;
    SS3[42][20] = 4'h0;
    SS3[43][20] = 4'h0;
    SS3[44][20] = 4'h0;
    SS3[45][20] = 4'h0;
    SS3[46][20] = 4'h0;
    SS3[47][20] = 4'h0;
    SS3[0][21] = 4'h0;
    SS3[1][21] = 4'hD;
    SS3[2][21] = 4'hD;
    SS3[3][21] = 4'hD;
    SS3[4][21] = 4'hC;
    SS3[5][21] = 4'hC;
    SS3[6][21] = 4'hC;
    SS3[7][21] = 4'hD;
    SS3[8][21] = 4'hD;
    SS3[9][21] = 4'hD;
    SS3[10][21] = 4'hC;
    SS3[11][21] = 4'hC;
    SS3[12][21] = 4'hC;
    SS3[13][21] = 4'hC;
    SS3[14][21] = 4'hC;
    SS3[15][21] = 4'hC;
    SS3[16][21] = 4'hC;
    SS3[17][21] = 4'hC;
    SS3[18][21] = 4'hC;
    SS3[19][21] = 4'hC;
    SS3[20][21] = 4'hC;
    SS3[21][21] = 4'hC;
    SS3[22][21] = 4'hC;
    SS3[23][21] = 4'hD;
    SS3[24][21] = 4'hD;
    SS3[25][21] = 4'hD;
    SS3[26][21] = 4'hA;
    SS3[27][21] = 4'hA;
    SS3[28][21] = 4'hA;
    SS3[29][21] = 4'hC;
    SS3[30][21] = 4'hC;
    SS3[31][21] = 4'hC;
    SS3[32][21] = 4'hC;
    SS3[33][21] = 4'hC;
    SS3[34][21] = 4'hC;
    SS3[35][21] = 4'hC;
    SS3[36][21] = 4'hC;
    SS3[37][21] = 4'hC;
    SS3[38][21] = 4'hD;
    SS3[39][21] = 4'hD;
    SS3[40][21] = 4'hD;
    SS3[41][21] = 4'hD;
    SS3[42][21] = 4'h0;
    SS3[43][21] = 4'h0;
    SS3[44][21] = 4'h0;
    SS3[45][21] = 4'h0;
    SS3[46][21] = 4'h0;
    SS3[47][21] = 4'h0;
    SS3[0][22] = 4'h0;
    SS3[1][22] = 4'hD;
    SS3[2][22] = 4'hD;
    SS3[3][22] = 4'hD;
    SS3[4][22] = 4'hE;
    SS3[5][22] = 4'hE;
    SS3[6][22] = 4'hE;
    SS3[7][22] = 4'hD;
    SS3[8][22] = 4'hD;
    SS3[9][22] = 4'hD;
    SS3[10][22] = 4'hD;
    SS3[11][22] = 4'hC;
    SS3[12][22] = 4'hD;
    SS3[13][22] = 4'hD;
    SS3[14][22] = 4'hC;
    SS3[15][22] = 4'hC;
    SS3[16][22] = 4'hC;
    SS3[17][22] = 4'hC;
    SS3[18][22] = 4'hC;
    SS3[19][22] = 4'hC;
    SS3[20][22] = 4'hC;
    SS3[21][22] = 4'hC;
    SS3[22][22] = 4'hC;
    SS3[23][22] = 4'hD;
    SS3[24][22] = 4'hD;
    SS3[25][22] = 4'hD;
    SS3[26][22] = 4'hD;
    SS3[27][22] = 4'hA;
    SS3[28][22] = 4'hA;
    SS3[29][22] = 4'hA;
    SS3[30][22] = 4'hC;
    SS3[31][22] = 4'hC;
    SS3[32][22] = 4'hC;
    SS3[33][22] = 4'hC;
    SS3[34][22] = 4'hC;
    SS3[35][22] = 4'hD;
    SS3[36][22] = 4'hD;
    SS3[37][22] = 4'hD;
    SS3[38][22] = 4'hD;
    SS3[39][22] = 4'hD;
    SS3[40][22] = 4'hD;
    SS3[41][22] = 4'hD;
    SS3[42][22] = 4'hD;
    SS3[43][22] = 4'h0;
    SS3[44][22] = 4'h0;
    SS3[45][22] = 4'h0;
    SS3[46][22] = 4'h0;
    SS3[47][22] = 4'h0;
    SS3[0][23] = 4'h0;
    SS3[1][23] = 4'hD;
    SS3[2][23] = 4'h0;
    SS3[3][23] = 4'h0;
    SS3[4][23] = 4'h0;
    SS3[5][23] = 4'hE;
    SS3[6][23] = 4'hE;
    SS3[7][23] = 4'hE;
    SS3[8][23] = 4'hD;
    SS3[9][23] = 4'hD;
    SS3[10][23] = 4'hE;
    SS3[11][23] = 4'hD;
    SS3[12][23] = 4'hD;
    SS3[13][23] = 4'hD;
    SS3[14][23] = 4'hC;
    SS3[15][23] = 4'hC;
    SS3[16][23] = 4'hC;
    SS3[17][23] = 4'hD;
    SS3[18][23] = 4'hD;
    SS3[19][23] = 4'hD;
    SS3[20][23] = 4'hD;
    SS3[21][23] = 4'hC;
    SS3[22][23] = 4'hC;
    SS3[23][23] = 4'hC;
    SS3[24][23] = 4'hD;
    SS3[25][23] = 4'hD;
    SS3[26][23] = 4'hD;
    SS3[27][23] = 4'hA;
    SS3[28][23] = 4'hA;
    SS3[29][23] = 4'hA;
    SS3[30][23] = 4'hC;
    SS3[31][23] = 4'hC;
    SS3[32][23] = 4'hC;
    SS3[33][23] = 4'hD;
    SS3[34][23] = 4'hD;
    SS3[35][23] = 4'hD;
    SS3[36][23] = 4'hD;
    SS3[37][23] = 4'hD;
    SS3[38][23] = 4'hD;
    SS3[39][23] = 4'hD;
    SS3[40][23] = 4'hD;
    SS3[41][23] = 4'h0;
    SS3[42][23] = 4'h0;
    SS3[43][23] = 4'h0;
    SS3[44][23] = 4'h0;
    SS3[45][23] = 4'h0;
    SS3[46][23] = 4'h0;
    SS3[47][23] = 4'h0;
    SS3[0][24] = 4'h0;
    SS3[1][24] = 4'h0;
    SS3[2][24] = 4'h0;
    SS3[3][24] = 4'h0;
    SS3[4][24] = 4'h0;
    SS3[5][24] = 4'hE;
    SS3[6][24] = 4'hE;
    SS3[7][24] = 4'h0;
    SS3[8][24] = 4'hE;
    SS3[9][24] = 4'hE;
    SS3[10][24] = 4'hE;
    SS3[11][24] = 4'hD;
    SS3[12][24] = 4'hD;
    SS3[13][24] = 4'hD;
    SS3[14][24] = 4'hD;
    SS3[15][24] = 4'hE;
    SS3[16][24] = 4'hE;
    SS3[17][24] = 4'hE;
    SS3[18][24] = 4'hD;
    SS3[19][24] = 4'hD;
    SS3[20][24] = 4'hD;
    SS3[21][24] = 4'hC;
    SS3[22][24] = 4'hC;
    SS3[23][24] = 4'hC;
    SS3[24][24] = 4'hD;
    SS3[25][24] = 4'hD;
    SS3[26][24] = 4'hD;
    SS3[27][24] = 4'hA;
    SS3[28][24] = 4'hA;
    SS3[29][24] = 4'hA;
    SS3[30][24] = 4'hA;
    SS3[31][24] = 4'hC;
    SS3[32][24] = 4'hC;
    SS3[33][24] = 4'hC;
    SS3[34][24] = 4'hD;
    SS3[35][24] = 4'hD;
    SS3[36][24] = 4'hD;
    SS3[37][24] = 4'hD;
    SS3[38][24] = 4'h0;
    SS3[39][24] = 4'h0;
    SS3[40][24] = 4'h0;
    SS3[41][24] = 4'h0;
    SS3[42][24] = 4'h0;
    SS3[43][24] = 4'h0;
    SS3[44][24] = 4'h0;
    SS3[45][24] = 4'h0;
    SS3[46][24] = 4'h0;
    SS3[47][24] = 4'h0;
    SS3[0][25] = 4'h0;
    SS3[1][25] = 4'h0;
    SS3[2][25] = 4'h0;
    SS3[3][25] = 4'h0;
    SS3[4][25] = 4'h0;
    SS3[5][25] = 4'h0;
    SS3[6][25] = 4'h0;
    SS3[7][25] = 4'h0;
    SS3[8][25] = 4'h0;
    SS3[9][25] = 4'hE;
    SS3[10][25] = 4'hE;
    SS3[11][25] = 4'hE;
    SS3[12][25] = 4'hD;
    SS3[13][25] = 4'hE;
    SS3[14][25] = 4'hE;
    SS3[15][25] = 4'hE;
    SS3[16][25] = 4'hE;
    SS3[17][25] = 4'hE;
    SS3[18][25] = 4'hD;
    SS3[19][25] = 4'hD;
    SS3[20][25] = 4'hD;
    SS3[21][25] = 4'hC;
    SS3[22][25] = 4'hC;
    SS3[23][25] = 4'hC;
    SS3[24][25] = 4'hC;
    SS3[25][25] = 4'hD;
    SS3[26][25] = 4'hD;
    SS3[27][25] = 4'hD;
    SS3[28][25] = 4'hD;
    SS3[29][25] = 4'hD;
    SS3[30][25] = 4'hD;
    SS3[31][25] = 4'hC;
    SS3[32][25] = 4'hC;
    SS3[33][25] = 4'hC;
    SS3[34][25] = 4'hD;
    SS3[35][25] = 4'hD;
    SS3[36][25] = 4'h0;
    SS3[37][25] = 4'h0;
    SS3[38][25] = 4'h0;
    SS3[39][25] = 4'h0;
    SS3[40][25] = 4'h0;
    SS3[41][25] = 4'h0;
    SS3[42][25] = 4'h0;
    SS3[43][25] = 4'h0;
    SS3[44][25] = 4'h0;
    SS3[45][25] = 4'h0;
    SS3[46][25] = 4'h0;
    SS3[47][25] = 4'h0;
    SS3[0][26] = 4'h0;
    SS3[1][26] = 4'h0;
    SS3[2][26] = 4'h0;
    SS3[3][26] = 4'h0;
    SS3[4][26] = 4'h0;
    SS3[5][26] = 4'h0;
    SS3[6][26] = 4'h0;
    SS3[7][26] = 4'h0;
    SS3[8][26] = 4'h0;
    SS3[9][26] = 4'hE;
    SS3[10][26] = 4'h0;
    SS3[11][26] = 4'h0;
    SS3[12][26] = 4'hE;
    SS3[13][26] = 4'hE;
    SS3[14][26] = 4'hE;
    SS3[15][26] = 4'hE;
    SS3[16][26] = 4'hE;
    SS3[17][26] = 4'hE;
    SS3[18][26] = 4'hE;
    SS3[19][26] = 4'hD;
    SS3[20][26] = 4'hD;
    SS3[21][26] = 4'hD;
    SS3[22][26] = 4'hC;
    SS3[23][26] = 4'hC;
    SS3[24][26] = 4'hC;
    SS3[25][26] = 4'hD;
    SS3[26][26] = 4'hC;
    SS3[27][26] = 4'hC;
    SS3[28][26] = 4'hD;
    SS3[29][26] = 4'hD;
    SS3[30][26] = 4'hD;
    SS3[31][26] = 4'hC;
    SS3[32][26] = 4'hC;
    SS3[33][26] = 4'hE;
    SS3[34][26] = 4'h0;
    SS3[35][26] = 4'h0;
    SS3[36][26] = 4'h0;
    SS3[37][26] = 4'h0;
    SS3[38][26] = 4'h0;
    SS3[39][26] = 4'h0;
    SS3[40][26] = 4'h0;
    SS3[41][26] = 4'h0;
    SS3[42][26] = 4'h0;
    SS3[43][26] = 4'h0;
    SS3[44][26] = 4'h0;
    SS3[45][26] = 4'h0;
    SS3[46][26] = 4'h0;
    SS3[47][26] = 4'h0;
    SS3[0][27] = 4'h0;
    SS3[1][27] = 4'h0;
    SS3[2][27] = 4'h0;
    SS3[3][27] = 4'h0;
    SS3[4][27] = 4'h0;
    SS3[5][27] = 4'h0;
    SS3[6][27] = 4'h0;
    SS3[7][27] = 4'h0;
    SS3[8][27] = 4'h0;
    SS3[9][27] = 4'h0;
    SS3[10][27] = 4'h0;
    SS3[11][27] = 4'h0;
    SS3[12][27] = 4'h0;
    SS3[13][27] = 4'hE;
    SS3[14][27] = 4'hE;
    SS3[15][27] = 4'hE;
    SS3[16][27] = 4'hE;
    SS3[17][27] = 4'hE;
    SS3[18][27] = 4'hE;
    SS3[19][27] = 4'hD;
    SS3[20][27] = 4'hD;
    SS3[21][27] = 4'hD;
    SS3[22][27] = 4'hC;
    SS3[23][27] = 4'hC;
    SS3[24][27] = 4'hC;
    SS3[25][27] = 4'hC;
    SS3[26][27] = 4'hC;
    SS3[27][27] = 4'hC;
    SS3[28][27] = 4'hC;
    SS3[29][27] = 4'hD;
    SS3[30][27] = 4'hD;
    SS3[31][27] = 4'hD;
    SS3[32][27] = 4'h0;
    SS3[33][27] = 4'h0;
    SS3[34][27] = 4'h0;
    SS3[35][27] = 4'h0;
    SS3[36][27] = 4'h0;
    SS3[37][27] = 4'h0;
    SS3[38][27] = 4'h0;
    SS3[39][27] = 4'h0;
    SS3[40][27] = 4'h0;
    SS3[41][27] = 4'h0;
    SS3[42][27] = 4'h0;
    SS3[43][27] = 4'h0;
    SS3[44][27] = 4'h0;
    SS3[45][27] = 4'h0;
    SS3[46][27] = 4'h0;
    SS3[47][27] = 4'h0;
    SS3[0][28] = 4'h0;
    SS3[1][28] = 4'h0;
    SS3[2][28] = 4'h0;
    SS3[3][28] = 4'h0;
    SS3[4][28] = 4'h0;
    SS3[5][28] = 4'h0;
    SS3[6][28] = 4'h0;
    SS3[7][28] = 4'h0;
    SS3[8][28] = 4'h0;
    SS3[9][28] = 4'h0;
    SS3[10][28] = 4'h0;
    SS3[11][28] = 4'h0;
    SS3[12][28] = 4'h0;
    SS3[13][28] = 4'hE;
    SS3[14][28] = 4'hE;
    SS3[15][28] = 4'hE;
    SS3[16][28] = 4'hE;
    SS3[17][28] = 4'hE;
    SS3[18][28] = 4'hE;
    SS3[19][28] = 4'hD;
    SS3[20][28] = 4'hD;
    SS3[21][28] = 4'hC;
    SS3[22][28] = 4'hC;
    SS3[23][28] = 4'hC;
    SS3[24][28] = 4'hC;
    SS3[25][28] = 4'hC;
    SS3[26][28] = 4'hC;
    SS3[27][28] = 4'hC;
    SS3[28][28] = 4'hC;
    SS3[29][28] = 4'hD;
    SS3[30][28] = 4'hD;
    SS3[31][28] = 4'hD;
    SS3[32][28] = 4'h0;
    SS3[33][28] = 4'h0;
    SS3[34][28] = 4'h0;
    SS3[35][28] = 4'h0;
    SS3[36][28] = 4'h0;
    SS3[37][28] = 4'h0;
    SS3[38][28] = 4'h0;
    SS3[39][28] = 4'h0;
    SS3[40][28] = 4'h0;
    SS3[41][28] = 4'h0;
    SS3[42][28] = 4'h0;
    SS3[43][28] = 4'h0;
    SS3[44][28] = 4'h0;
    SS3[45][28] = 4'h0;
    SS3[46][28] = 4'h0;
    SS3[47][28] = 4'h0;
    SS3[0][29] = 4'h0;
    SS3[1][29] = 4'h0;
    SS3[2][29] = 4'h0;
    SS3[3][29] = 4'h0;
    SS3[4][29] = 4'h0;
    SS3[5][29] = 4'h0;
    SS3[6][29] = 4'h0;
    SS3[7][29] = 4'h0;
    SS3[8][29] = 4'h0;
    SS3[9][29] = 4'h0;
    SS3[10][29] = 4'h0;
    SS3[11][29] = 4'h0;
    SS3[12][29] = 4'h0;
    SS3[13][29] = 4'hE;
    SS3[14][29] = 4'hE;
    SS3[15][29] = 4'hE;
    SS3[16][29] = 4'hE;
    SS3[17][29] = 4'hE;
    SS3[18][29] = 4'hC;
    SS3[19][29] = 4'hC;
    SS3[20][29] = 4'hC;
    SS3[21][29] = 4'hC;
    SS3[22][29] = 4'hC;
    SS3[23][29] = 4'hC;
    SS3[24][29] = 4'hC;
    SS3[25][29] = 4'hC;
    SS3[26][29] = 4'hD;
    SS3[27][29] = 4'hD;
    SS3[28][29] = 4'hD;
    SS3[29][29] = 4'hD;
    SS3[30][29] = 4'hD;
    SS3[31][29] = 4'hD;
    SS3[32][29] = 4'hD;
    SS3[33][29] = 4'h0;
    SS3[34][29] = 4'h0;
    SS3[35][29] = 4'h0;
    SS3[36][29] = 4'h0;
    SS3[37][29] = 4'h0;
    SS3[38][29] = 4'h0;
    SS3[39][29] = 4'h0;
    SS3[40][29] = 4'h0;
    SS3[41][29] = 4'h0;
    SS3[42][29] = 4'h0;
    SS3[43][29] = 4'h0;
    SS3[44][29] = 4'h0;
    SS3[45][29] = 4'h0;
    SS3[46][29] = 4'h0;
    SS3[47][29] = 4'h0;
    SS3[0][30] = 4'h0;
    SS3[1][30] = 4'h0;
    SS3[2][30] = 4'h0;
    SS3[3][30] = 4'h0;
    SS3[4][30] = 4'h0;
    SS3[5][30] = 4'h0;
    SS3[6][30] = 4'h0;
    SS3[7][30] = 4'h0;
    SS3[8][30] = 4'h0;
    SS3[9][30] = 4'h0;
    SS3[10][30] = 4'h0;
    SS3[11][30] = 4'h0;
    SS3[12][30] = 4'h0;
    SS3[13][30] = 4'h0;
    SS3[14][30] = 4'hE;
    SS3[15][30] = 4'hE;
    SS3[16][30] = 4'hD;
    SS3[17][30] = 4'hC;
    SS3[18][30] = 4'hC;
    SS3[19][30] = 4'hC;
    SS3[20][30] = 4'hC;
    SS3[21][30] = 4'hC;
    SS3[22][30] = 4'hC;
    SS3[23][30] = 4'hC;
    SS3[24][30] = 4'hE;
    SS3[25][30] = 4'hE;
    SS3[26][30] = 4'hE;
    SS3[27][30] = 4'hD;
    SS3[28][30] = 4'hD;
    SS3[29][30] = 4'hD;
    SS3[30][30] = 4'hD;
    SS3[31][30] = 4'hD;
    SS3[32][30] = 4'h3;
    SS3[33][30] = 4'h0;
    SS3[34][30] = 4'h0;
    SS3[35][30] = 4'h0;
    SS3[36][30] = 4'h0;
    SS3[37][30] = 4'h0;
    SS3[38][30] = 4'h0;
    SS3[39][30] = 4'h0;
    SS3[40][30] = 4'h0;
    SS3[41][30] = 4'h0;
    SS3[42][30] = 4'h0;
    SS3[43][30] = 4'h0;
    SS3[44][30] = 4'h0;
    SS3[45][30] = 4'h0;
    SS3[46][30] = 4'h0;
    SS3[47][30] = 4'h0;
    SS3[0][31] = 4'h0;
    SS3[1][31] = 4'h0;
    SS3[2][31] = 4'h0;
    SS3[3][31] = 4'h0;
    SS3[4][31] = 4'h0;
    SS3[5][31] = 4'h0;
    SS3[6][31] = 4'h0;
    SS3[7][31] = 4'h0;
    SS3[8][31] = 4'h0;
    SS3[9][31] = 4'h0;
    SS3[10][31] = 4'h0;
    SS3[11][31] = 4'h0;
    SS3[12][31] = 4'h0;
    SS3[13][31] = 4'h0;
    SS3[14][31] = 4'hD;
    SS3[15][31] = 4'hD;
    SS3[16][31] = 4'hD;
    SS3[17][31] = 4'hC;
    SS3[18][31] = 4'hC;
    SS3[19][31] = 4'hC;
    SS3[20][31] = 4'hC;
    SS3[21][31] = 4'hC;
    SS3[22][31] = 4'hC;
    SS3[23][31] = 4'hC;
    SS3[24][31] = 4'hE;
    SS3[25][31] = 4'hE;
    SS3[26][31] = 4'hE;
    SS3[27][31] = 4'hD;
    SS3[28][31] = 4'hD;
    SS3[29][31] = 4'hD;
    SS3[30][31] = 4'h3;
    SS3[31][31] = 4'h3;
    SS3[32][31] = 4'h3;
    SS3[33][31] = 4'h3;
    SS3[34][31] = 4'h0;
    SS3[35][31] = 4'h0;
    SS3[36][31] = 4'h0;
    SS3[37][31] = 4'h0;
    SS3[38][31] = 4'h0;
    SS3[39][31] = 4'h0;
    SS3[40][31] = 4'h0;
    SS3[41][31] = 4'h0;
    SS3[42][31] = 4'h0;
    SS3[43][31] = 4'h0;
    SS3[44][31] = 4'h0;
    SS3[45][31] = 4'h0;
    SS3[46][31] = 4'h0;
    SS3[47][31] = 4'h0;
    SS3[0][32] = 4'h0;
    SS3[1][32] = 4'h0;
    SS3[2][32] = 4'h0;
    SS3[3][32] = 4'h0;
    SS3[4][32] = 4'h0;
    SS3[5][32] = 4'h0;
    SS3[6][32] = 4'h0;
    SS3[7][32] = 4'h0;
    SS3[8][32] = 4'h0;
    SS3[9][32] = 4'h0;
    SS3[10][32] = 4'h0;
    SS3[11][32] = 4'hE;
    SS3[12][32] = 4'hE;
    SS3[13][32] = 4'hE;
    SS3[14][32] = 4'hE;
    SS3[15][32] = 4'hD;
    SS3[16][32] = 4'hD;
    SS3[17][32] = 4'hD;
    SS3[18][32] = 4'hC;
    SS3[19][32] = 4'hC;
    SS3[20][32] = 4'hC;
    SS3[21][32] = 4'hC;
    SS3[22][32] = 4'hC;
    SS3[23][32] = 4'hC;
    SS3[24][32] = 4'hE;
    SS3[25][32] = 4'hE;
    SS3[26][32] = 4'hE;
    SS3[27][32] = 4'hD;
    SS3[28][32] = 4'hD;
    SS3[29][32] = 4'hD;
    SS3[30][32] = 4'hD;
    SS3[31][32] = 4'h3;
    SS3[32][32] = 4'h3;
    SS3[33][32] = 4'h3;
    SS3[34][32] = 4'h0;
    SS3[35][32] = 4'h0;
    SS3[36][32] = 4'h0;
    SS3[37][32] = 4'h0;
    SS3[38][32] = 4'h0;
    SS3[39][32] = 4'h0;
    SS3[40][32] = 4'h0;
    SS3[41][32] = 4'h0;
    SS3[42][32] = 4'h0;
    SS3[43][32] = 4'h0;
    SS3[44][32] = 4'h0;
    SS3[45][32] = 4'h0;
    SS3[46][32] = 4'h0;
    SS3[47][32] = 4'h0;
    SS3[0][33] = 4'h0;
    SS3[1][33] = 4'h0;
    SS3[2][33] = 4'h0;
    SS3[3][33] = 4'h0;
    SS3[4][33] = 4'h0;
    SS3[5][33] = 4'h0;
    SS3[6][33] = 4'h0;
    SS3[7][33] = 4'h0;
    SS3[8][33] = 4'h0;
    SS3[9][33] = 4'h0;
    SS3[10][33] = 4'h0;
    SS3[11][33] = 4'h0;
    SS3[12][33] = 4'hE;
    SS3[13][33] = 4'hE;
    SS3[14][33] = 4'hE;
    SS3[15][33] = 4'hD;
    SS3[16][33] = 4'hD;
    SS3[17][33] = 4'hC;
    SS3[18][33] = 4'hC;
    SS3[19][33] = 4'hC;
    SS3[20][33] = 4'hC;
    SS3[21][33] = 4'hC;
    SS3[22][33] = 4'hC;
    SS3[23][33] = 4'hC;
    SS3[24][33] = 4'hE;
    SS3[25][33] = 4'hD;
    SS3[26][33] = 4'hD;
    SS3[27][33] = 4'hD;
    SS3[28][33] = 4'hD;
    SS3[29][33] = 4'hD;
    SS3[30][33] = 4'hD;
    SS3[31][33] = 4'h3;
    SS3[32][33] = 4'h0;
    SS3[33][33] = 4'h0;
    SS3[34][33] = 4'h0;
    SS3[35][33] = 4'h0;
    SS3[36][33] = 4'h0;
    SS3[37][33] = 4'h0;
    SS3[38][33] = 4'h0;
    SS3[39][33] = 4'h0;
    SS3[40][33] = 4'h0;
    SS3[41][33] = 4'h0;
    SS3[42][33] = 4'h0;
    SS3[43][33] = 4'h0;
    SS3[44][33] = 4'h0;
    SS3[45][33] = 4'h0;
    SS3[46][33] = 4'h0;
    SS3[47][33] = 4'h0;
    SS3[0][34] = 4'h0;
    SS3[1][34] = 4'h0;
    SS3[2][34] = 4'h0;
    SS3[3][34] = 4'h0;
    SS3[4][34] = 4'h0;
    SS3[5][34] = 4'h0;
    SS3[6][34] = 4'h0;
    SS3[7][34] = 4'h0;
    SS3[8][34] = 4'h0;
    SS3[9][34] = 4'h0;
    SS3[10][34] = 4'h0;
    SS3[11][34] = 4'h0;
    SS3[12][34] = 4'hE;
    SS3[13][34] = 4'hE;
    SS3[14][34] = 4'hD;
    SS3[15][34] = 4'hD;
    SS3[16][34] = 4'hC;
    SS3[17][34] = 4'hC;
    SS3[18][34] = 4'hC;
    SS3[19][34] = 4'hC;
    SS3[20][34] = 4'hC;
    SS3[21][34] = 4'hC;
    SS3[22][34] = 4'hE;
    SS3[23][34] = 4'hE;
    SS3[24][34] = 4'hE;
    SS3[25][34] = 4'hD;
    SS3[26][34] = 4'hD;
    SS3[27][34] = 4'hD;
    SS3[28][34] = 4'hD;
    SS3[29][34] = 4'hD;
    SS3[30][34] = 4'h0;
    SS3[31][34] = 4'h0;
    SS3[32][34] = 4'h0;
    SS3[33][34] = 4'h0;
    SS3[34][34] = 4'h0;
    SS3[35][34] = 4'h0;
    SS3[36][34] = 4'h0;
    SS3[37][34] = 4'h0;
    SS3[38][34] = 4'h0;
    SS3[39][34] = 4'h0;
    SS3[40][34] = 4'h0;
    SS3[41][34] = 4'h0;
    SS3[42][34] = 4'h0;
    SS3[43][34] = 4'h0;
    SS3[44][34] = 4'h0;
    SS3[45][34] = 4'h0;
    SS3[46][34] = 4'h0;
    SS3[47][34] = 4'h0;
    SS3[0][35] = 4'h0;
    SS3[1][35] = 4'h0;
    SS3[2][35] = 4'h0;
    SS3[3][35] = 4'h0;
    SS3[4][35] = 4'h0;
    SS3[5][35] = 4'h0;
    SS3[6][35] = 4'h0;
    SS3[7][35] = 4'h0;
    SS3[8][35] = 4'h0;
    SS3[9][35] = 4'h0;
    SS3[10][35] = 4'h0;
    SS3[11][35] = 4'h0;
    SS3[12][35] = 4'hE;
    SS3[13][35] = 4'hD;
    SS3[14][35] = 4'hD;
    SS3[15][35] = 4'hD;
    SS3[16][35] = 4'hC;
    SS3[17][35] = 4'hC;
    SS3[18][35] = 4'hC;
    SS3[19][35] = 4'hC;
    SS3[20][35] = 4'hC;
    SS3[21][35] = 4'hC;
    SS3[22][35] = 4'hE;
    SS3[23][35] = 4'hE;
    SS3[24][35] = 4'hE;
    SS3[25][35] = 4'hE;
    SS3[26][35] = 4'hD;
    SS3[27][35] = 4'hD;
    SS3[28][35] = 4'hD;
    SS3[29][35] = 4'h0;
    SS3[30][35] = 4'h0;
    SS3[31][35] = 4'h0;
    SS3[32][35] = 4'h0;
    SS3[33][35] = 4'h0;
    SS3[34][35] = 4'h0;
    SS3[35][35] = 4'h0;
    SS3[36][35] = 4'h0;
    SS3[37][35] = 4'h0;
    SS3[38][35] = 4'h0;
    SS3[39][35] = 4'h0;
    SS3[40][35] = 4'h0;
    SS3[41][35] = 4'h0;
    SS3[42][35] = 4'h0;
    SS3[43][35] = 4'h0;
    SS3[44][35] = 4'h0;
    SS3[45][35] = 4'h0;
    SS3[46][35] = 4'h0;
    SS3[47][35] = 4'h0;
    SS3[0][36] = 4'h0;
    SS3[1][36] = 4'h0;
    SS3[2][36] = 4'h0;
    SS3[3][36] = 4'h0;
    SS3[4][36] = 4'h0;
    SS3[5][36] = 4'h0;
    SS3[6][36] = 4'h0;
    SS3[7][36] = 4'h0;
    SS3[8][36] = 4'h0;
    SS3[9][36] = 4'h0;
    SS3[10][36] = 4'hE;
    SS3[11][36] = 4'hE;
    SS3[12][36] = 4'hE;
    SS3[13][36] = 4'hD;
    SS3[14][36] = 4'hD;
    SS3[15][36] = 4'hD;
    SS3[16][36] = 4'hC;
    SS3[17][36] = 4'hC;
    SS3[18][36] = 4'hC;
    SS3[19][36] = 4'hC;
    SS3[20][36] = 4'hC;
    SS3[21][36] = 4'hC;
    SS3[22][36] = 4'hC;
    SS3[23][36] = 4'hE;
    SS3[24][36] = 4'hE;
    SS3[25][36] = 4'hE;
    SS3[26][36] = 4'hD;
    SS3[27][36] = 4'hD;
    SS3[28][36] = 4'hD;
    SS3[29][36] = 4'h0;
    SS3[30][36] = 4'h0;
    SS3[31][36] = 4'h0;
    SS3[32][36] = 4'h0;
    SS3[33][36] = 4'h0;
    SS3[34][36] = 4'h0;
    SS3[35][36] = 4'h0;
    SS3[36][36] = 4'h0;
    SS3[37][36] = 4'h0;
    SS3[38][36] = 4'h0;
    SS3[39][36] = 4'h0;
    SS3[40][36] = 4'h0;
    SS3[41][36] = 4'h0;
    SS3[42][36] = 4'h0;
    SS3[43][36] = 4'h0;
    SS3[44][36] = 4'h0;
    SS3[45][36] = 4'h0;
    SS3[46][36] = 4'h0;
    SS3[47][36] = 4'h0;
    SS3[0][37] = 4'h0;
    SS3[1][37] = 4'h0;
    SS3[2][37] = 4'h0;
    SS3[3][37] = 4'h0;
    SS3[4][37] = 4'h0;
    SS3[5][37] = 4'h0;
    SS3[6][37] = 4'h0;
    SS3[7][37] = 4'h0;
    SS3[8][37] = 4'h0;
    SS3[9][37] = 4'h0;
    SS3[10][37] = 4'hE;
    SS3[11][37] = 4'hE;
    SS3[12][37] = 4'hE;
    SS3[13][37] = 4'hE;
    SS3[14][37] = 4'hD;
    SS3[15][37] = 4'hC;
    SS3[16][37] = 4'hC;
    SS3[17][37] = 4'hC;
    SS3[18][37] = 4'hC;
    SS3[19][37] = 4'hC;
    SS3[20][37] = 4'hC;
    SS3[21][37] = 4'hC;
    SS3[22][37] = 4'hE;
    SS3[23][37] = 4'hE;
    SS3[24][37] = 4'hE;
    SS3[25][37] = 4'hE;
    SS3[26][37] = 4'hD;
    SS3[27][37] = 4'hD;
    SS3[28][37] = 4'hD;
    SS3[29][37] = 4'hD;
    SS3[30][37] = 4'h0;
    SS3[31][37] = 4'h0;
    SS3[32][37] = 4'h0;
    SS3[33][37] = 4'h0;
    SS3[34][37] = 4'h0;
    SS3[35][37] = 4'h0;
    SS3[36][37] = 4'h0;
    SS3[37][37] = 4'h0;
    SS3[38][37] = 4'h0;
    SS3[39][37] = 4'h0;
    SS3[40][37] = 4'h0;
    SS3[41][37] = 4'h0;
    SS3[42][37] = 4'h0;
    SS3[43][37] = 4'h0;
    SS3[44][37] = 4'h0;
    SS3[45][37] = 4'h0;
    SS3[46][37] = 4'h0;
    SS3[47][37] = 4'h0;
    SS3[0][38] = 4'h0;
    SS3[1][38] = 4'h0;
    SS3[2][38] = 4'h0;
    SS3[3][38] = 4'h0;
    SS3[4][38] = 4'h0;
    SS3[5][38] = 4'h0;
    SS3[6][38] = 4'h0;
    SS3[7][38] = 4'h0;
    SS3[8][38] = 4'h0;
    SS3[9][38] = 4'h0;
    SS3[10][38] = 4'h0;
    SS3[11][38] = 4'hE;
    SS3[12][38] = 4'hC;
    SS3[13][38] = 4'hC;
    SS3[14][38] = 4'hC;
    SS3[15][38] = 4'hC;
    SS3[16][38] = 4'hC;
    SS3[17][38] = 4'hC;
    SS3[18][38] = 4'hC;
    SS3[19][38] = 4'hC;
    SS3[20][38] = 4'hE;
    SS3[21][38] = 4'hE;
    SS3[22][38] = 4'hE;
    SS3[23][38] = 4'hE;
    SS3[24][38] = 4'hE;
    SS3[25][38] = 4'hE;
    SS3[26][38] = 4'hE;
    SS3[27][38] = 4'hD;
    SS3[28][38] = 4'h3;
    SS3[29][38] = 4'h3;
    SS3[30][38] = 4'h0;
    SS3[31][38] = 4'h0;
    SS3[32][38] = 4'h0;
    SS3[33][38] = 4'h0;
    SS3[34][38] = 4'h0;
    SS3[35][38] = 4'h0;
    SS3[36][38] = 4'h0;
    SS3[37][38] = 4'h0;
    SS3[38][38] = 4'h0;
    SS3[39][38] = 4'h0;
    SS3[40][38] = 4'h0;
    SS3[41][38] = 4'h0;
    SS3[42][38] = 4'h0;
    SS3[43][38] = 4'h0;
    SS3[44][38] = 4'h0;
    SS3[45][38] = 4'h0;
    SS3[46][38] = 4'h0;
    SS3[47][38] = 4'h0;
    SS3[0][39] = 4'h0;
    SS3[1][39] = 4'h0;
    SS3[2][39] = 4'h0;
    SS3[3][39] = 4'h0;
    SS3[4][39] = 4'h0;
    SS3[5][39] = 4'h0;
    SS3[6][39] = 4'h0;
    SS3[7][39] = 4'h0;
    SS3[8][39] = 4'h0;
    SS3[9][39] = 4'h0;
    SS3[10][39] = 4'hD;
    SS3[11][39] = 4'hC;
    SS3[12][39] = 4'hC;
    SS3[13][39] = 4'hC;
    SS3[14][39] = 4'hC;
    SS3[15][39] = 4'hC;
    SS3[16][39] = 4'hC;
    SS3[17][39] = 4'hC;
    SS3[18][39] = 4'h0;
    SS3[19][39] = 4'h0;
    SS3[20][39] = 4'h0;
    SS3[21][39] = 4'hE;
    SS3[22][39] = 4'hE;
    SS3[23][39] = 4'hE;
    SS3[24][39] = 4'hE;
    SS3[25][39] = 4'hD;
    SS3[26][39] = 4'hD;
    SS3[27][39] = 4'h3;
    SS3[28][39] = 4'h3;
    SS3[29][39] = 4'h3;
    SS3[30][39] = 4'h0;
    SS3[31][39] = 4'h0;
    SS3[32][39] = 4'h0;
    SS3[33][39] = 4'h0;
    SS3[34][39] = 4'h0;
    SS3[35][39] = 4'h0;
    SS3[36][39] = 4'h0;
    SS3[37][39] = 4'h0;
    SS3[38][39] = 4'h0;
    SS3[39][39] = 4'h0;
    SS3[40][39] = 4'h0;
    SS3[41][39] = 4'h0;
    SS3[42][39] = 4'h0;
    SS3[43][39] = 4'h0;
    SS3[44][39] = 4'h0;
    SS3[45][39] = 4'h0;
    SS3[46][39] = 4'h0;
    SS3[47][39] = 4'h0;
    SS3[0][40] = 4'h0;
    SS3[1][40] = 4'h0;
    SS3[2][40] = 4'h0;
    SS3[3][40] = 4'h0;
    SS3[4][40] = 4'h0;
    SS3[5][40] = 4'h0;
    SS3[6][40] = 4'h0;
    SS3[7][40] = 4'h0;
    SS3[8][40] = 4'hD;
    SS3[9][40] = 4'hD;
    SS3[10][40] = 4'hD;
    SS3[11][40] = 4'hD;
    SS3[12][40] = 4'hC;
    SS3[13][40] = 4'hC;
    SS3[14][40] = 4'hC;
    SS3[15][40] = 4'h0;
    SS3[16][40] = 4'h0;
    SS3[17][40] = 4'h0;
    SS3[18][40] = 4'h0;
    SS3[19][40] = 4'h0;
    SS3[20][40] = 4'h0;
    SS3[21][40] = 4'hE;
    SS3[22][40] = 4'hE;
    SS3[23][40] = 4'hE;
    SS3[24][40] = 4'hD;
    SS3[25][40] = 4'hD;
    SS3[26][40] = 4'hD;
    SS3[27][40] = 4'hD;
    SS3[28][40] = 4'h3;
    SS3[29][40] = 4'h3;
    SS3[30][40] = 4'h3;
    SS3[31][40] = 4'h0;
    SS3[32][40] = 4'h0;
    SS3[33][40] = 4'h0;
    SS3[34][40] = 4'h0;
    SS3[35][40] = 4'h0;
    SS3[36][40] = 4'h0;
    SS3[37][40] = 4'h0;
    SS3[38][40] = 4'h0;
    SS3[39][40] = 4'h0;
    SS3[40][40] = 4'h0;
    SS3[41][40] = 4'h0;
    SS3[42][40] = 4'h0;
    SS3[43][40] = 4'h0;
    SS3[44][40] = 4'h0;
    SS3[45][40] = 4'h0;
    SS3[46][40] = 4'h0;
    SS3[47][40] = 4'h0;
    SS3[0][41] = 4'h0;
    SS3[1][41] = 4'h0;
    SS3[2][41] = 4'h0;
    SS3[3][41] = 4'h0;
    SS3[4][41] = 4'h0;
    SS3[5][41] = 4'h0;
    SS3[6][41] = 4'h0;
    SS3[7][41] = 4'h0;
    SS3[8][41] = 4'h0;
    SS3[9][41] = 4'hD;
    SS3[10][41] = 4'hD;
    SS3[11][41] = 4'hD;
    SS3[12][41] = 4'hC;
    SS3[13][41] = 4'hC;
    SS3[14][41] = 4'hC;
    SS3[15][41] = 4'h0;
    SS3[16][41] = 4'h0;
    SS3[17][41] = 4'h0;
    SS3[18][41] = 4'h0;
    SS3[19][41] = 4'h0;
    SS3[20][41] = 4'h0;
    SS3[21][41] = 4'h0;
    SS3[22][41] = 4'hE;
    SS3[23][41] = 4'hE;
    SS3[24][41] = 4'hE;
    SS3[25][41] = 4'hD;
    SS3[26][41] = 4'hD;
    SS3[27][41] = 4'hD;
    SS3[28][41] = 4'h0;
    SS3[29][41] = 4'h0;
    SS3[30][41] = 4'h0;
    SS3[31][41] = 4'h0;
    SS3[32][41] = 4'h0;
    SS3[33][41] = 4'h0;
    SS3[34][41] = 4'h0;
    SS3[35][41] = 4'h0;
    SS3[36][41] = 4'h0;
    SS3[37][41] = 4'h0;
    SS3[38][41] = 4'h0;
    SS3[39][41] = 4'h0;
    SS3[40][41] = 4'h0;
    SS3[41][41] = 4'h0;
    SS3[42][41] = 4'h0;
    SS3[43][41] = 4'h0;
    SS3[44][41] = 4'h0;
    SS3[45][41] = 4'h0;
    SS3[46][41] = 4'h0;
    SS3[47][41] = 4'h0;
    SS3[0][42] = 4'h0;
    SS3[1][42] = 4'h0;
    SS3[2][42] = 4'h0;
    SS3[3][42] = 4'h0;
    SS3[4][42] = 4'h0;
    SS3[5][42] = 4'h0;
    SS3[6][42] = 4'h0;
    SS3[7][42] = 4'h0;
    SS3[8][42] = 4'h0;
    SS3[9][42] = 4'hD;
    SS3[10][42] = 4'hC;
    SS3[11][42] = 4'hC;
    SS3[12][42] = 4'hC;
    SS3[13][42] = 4'hC;
    SS3[14][42] = 4'hC;
    SS3[15][42] = 4'hC;
    SS3[16][42] = 4'h0;
    SS3[17][42] = 4'h0;
    SS3[18][42] = 4'h0;
    SS3[19][42] = 4'h0;
    SS3[20][42] = 4'h0;
    SS3[21][42] = 4'h0;
    SS3[22][42] = 4'hE;
    SS3[23][42] = 4'hE;
    SS3[24][42] = 4'hE;
    SS3[25][42] = 4'hD;
    SS3[26][42] = 4'hD;
    SS3[27][42] = 4'hD;
    SS3[28][42] = 4'h0;
    SS3[29][42] = 4'h0;
    SS3[30][42] = 4'h0;
    SS3[31][42] = 4'h0;
    SS3[32][42] = 4'h0;
    SS3[33][42] = 4'h0;
    SS3[34][42] = 4'h0;
    SS3[35][42] = 4'h0;
    SS3[36][42] = 4'h0;
    SS3[37][42] = 4'h0;
    SS3[38][42] = 4'h0;
    SS3[39][42] = 4'h0;
    SS3[40][42] = 4'h0;
    SS3[41][42] = 4'h0;
    SS3[42][42] = 4'h0;
    SS3[43][42] = 4'h0;
    SS3[44][42] = 4'h0;
    SS3[45][42] = 4'h0;
    SS3[46][42] = 4'h0;
    SS3[47][42] = 4'h0;
    SS3[0][43] = 4'h0;
    SS3[1][43] = 4'h0;
    SS3[2][43] = 4'h0;
    SS3[3][43] = 4'h0;
    SS3[4][43] = 4'h0;
    SS3[5][43] = 4'h0;
    SS3[6][43] = 4'h0;
    SS3[7][43] = 4'h0;
    SS3[8][43] = 4'hD;
    SS3[9][43] = 4'hD;
    SS3[10][43] = 4'hC;
    SS3[11][43] = 4'hC;
    SS3[12][43] = 4'hC;
    SS3[13][43] = 4'hC;
    SS3[14][43] = 4'hC;
    SS3[15][43] = 4'hC;
    SS3[16][43] = 4'h0;
    SS3[17][43] = 4'h0;
    SS3[18][43] = 4'h0;
    SS3[19][43] = 4'h0;
    SS3[20][43] = 4'h0;
    SS3[21][43] = 4'h0;
    SS3[22][43] = 4'hE;
    SS3[23][43] = 4'hD;
    SS3[24][43] = 4'hD;
    SS3[25][43] = 4'hD;
    SS3[26][43] = 4'hD;
    SS3[27][43] = 4'hD;
    SS3[28][43] = 4'hD;
    SS3[29][43] = 4'h0;
    SS3[30][43] = 4'h0;
    SS3[31][43] = 4'h0;
    SS3[32][43] = 4'h0;
    SS3[33][43] = 4'h0;
    SS3[34][43] = 4'h0;
    SS3[35][43] = 4'h0;
    SS3[36][43] = 4'h0;
    SS3[37][43] = 4'h0;
    SS3[38][43] = 4'h0;
    SS3[39][43] = 4'h0;
    SS3[40][43] = 4'h0;
    SS3[41][43] = 4'h0;
    SS3[42][43] = 4'h0;
    SS3[43][43] = 4'h0;
    SS3[44][43] = 4'h0;
    SS3[45][43] = 4'h0;
    SS3[46][43] = 4'h0;
    SS3[47][43] = 4'h0;
    SS3[0][44] = 4'h0;
    SS3[1][44] = 4'h0;
    SS3[2][44] = 4'h0;
    SS3[3][44] = 4'h0;
    SS3[4][44] = 4'h0;
    SS3[5][44] = 4'h0;
    SS3[6][44] = 4'h0;
    SS3[7][44] = 4'hD;
    SS3[8][44] = 4'hD;
    SS3[9][44] = 4'hD;
    SS3[10][44] = 4'hC;
    SS3[11][44] = 4'hC;
    SS3[12][44] = 4'hC;
    SS3[13][44] = 4'h0;
    SS3[14][44] = 4'h0;
    SS3[15][44] = 4'h0;
    SS3[16][44] = 4'h0;
    SS3[17][44] = 4'h0;
    SS3[18][44] = 4'h0;
    SS3[19][44] = 4'h0;
    SS3[20][44] = 4'h0;
    SS3[21][44] = 4'h0;
    SS3[22][44] = 4'h0;
    SS3[23][44] = 4'hD;
    SS3[24][44] = 4'hD;
    SS3[25][44] = 4'hD;
    SS3[26][44] = 4'hD;
    SS3[27][44] = 4'hD;
    SS3[28][44] = 4'hD;
    SS3[29][44] = 4'h0;
    SS3[30][44] = 4'h0;
    SS3[31][44] = 4'h0;
    SS3[32][44] = 4'h0;
    SS3[33][44] = 4'h0;
    SS3[34][44] = 4'h0;
    SS3[35][44] = 4'h0;
    SS3[36][44] = 4'h0;
    SS3[37][44] = 4'h0;
    SS3[38][44] = 4'h0;
    SS3[39][44] = 4'h0;
    SS3[40][44] = 4'h0;
    SS3[41][44] = 4'h0;
    SS3[42][44] = 4'h0;
    SS3[43][44] = 4'h0;
    SS3[44][44] = 4'h0;
    SS3[45][44] = 4'h0;
    SS3[46][44] = 4'h0;
    SS3[47][44] = 4'h0;
    SS3[0][45] = 4'h0;
    SS3[1][45] = 4'h0;
    SS3[2][45] = 4'h0;
    SS3[3][45] = 4'h0;
    SS3[4][45] = 4'h0;
    SS3[5][45] = 4'h0;
    SS3[6][45] = 4'h0;
    SS3[7][45] = 4'hD;
    SS3[8][45] = 4'hD;
    SS3[9][45] = 4'hD;
    SS3[10][45] = 4'hC;
    SS3[11][45] = 4'h0;
    SS3[12][45] = 4'h0;
    SS3[13][45] = 4'h0;
    SS3[14][45] = 4'h0;
    SS3[15][45] = 4'h0;
    SS3[16][45] = 4'h0;
    SS3[17][45] = 4'h0;
    SS3[18][45] = 4'h0;
    SS3[19][45] = 4'h0;
    SS3[20][45] = 4'h0;
    SS3[21][45] = 4'h0;
    SS3[22][45] = 4'h0;
    SS3[23][45] = 4'hD;
    SS3[24][45] = 4'hD;
    SS3[25][45] = 4'hD;
    SS3[26][45] = 4'hE;
    SS3[27][45] = 4'h0;
    SS3[28][45] = 4'h0;
    SS3[29][45] = 4'h0;
    SS3[30][45] = 4'h0;
    SS3[31][45] = 4'h0;
    SS3[32][45] = 4'h0;
    SS3[33][45] = 4'h0;
    SS3[34][45] = 4'h0;
    SS3[35][45] = 4'h0;
    SS3[36][45] = 4'h0;
    SS3[37][45] = 4'h0;
    SS3[38][45] = 4'h0;
    SS3[39][45] = 4'h0;
    SS3[40][45] = 4'h0;
    SS3[41][45] = 4'h0;
    SS3[42][45] = 4'h0;
    SS3[43][45] = 4'h0;
    SS3[44][45] = 4'h0;
    SS3[45][45] = 4'h0;
    SS3[46][45] = 4'h0;
    SS3[47][45] = 4'h0;
    SS3[0][46] = 4'h0;
    SS3[1][46] = 4'h0;
    SS3[2][46] = 4'h0;
    SS3[3][46] = 4'h0;
    SS3[4][46] = 4'h0;
    SS3[5][46] = 4'h0;
    SS3[6][46] = 4'h0;
    SS3[7][46] = 4'h0;
    SS3[8][46] = 4'h0;
    SS3[9][46] = 4'h0;
    SS3[10][46] = 4'h0;
    SS3[11][46] = 4'h0;
    SS3[12][46] = 4'h0;
    SS3[13][46] = 4'h0;
    SS3[14][46] = 4'h0;
    SS3[15][46] = 4'h0;
    SS3[16][46] = 4'h0;
    SS3[17][46] = 4'h0;
    SS3[18][46] = 4'h0;
    SS3[19][46] = 4'h0;
    SS3[20][46] = 4'h0;
    SS3[21][46] = 4'h0;
    SS3[22][46] = 4'h0;
    SS3[23][46] = 4'h0;
    SS3[24][46] = 4'hD;
    SS3[25][46] = 4'hD;
    SS3[26][46] = 4'hD;
    SS3[27][46] = 4'h0;
    SS3[28][46] = 4'h0;
    SS3[29][46] = 4'h0;
    SS3[30][46] = 4'h0;
    SS3[31][46] = 4'h0;
    SS3[32][46] = 4'h0;
    SS3[33][46] = 4'h0;
    SS3[34][46] = 4'h0;
    SS3[35][46] = 4'h0;
    SS3[36][46] = 4'h0;
    SS3[37][46] = 4'h0;
    SS3[38][46] = 4'h0;
    SS3[39][46] = 4'h0;
    SS3[40][46] = 4'h0;
    SS3[41][46] = 4'h0;
    SS3[42][46] = 4'h0;
    SS3[43][46] = 4'h0;
    SS3[44][46] = 4'h0;
    SS3[45][46] = 4'h0;
    SS3[46][46] = 4'h0;
    SS3[47][46] = 4'h0;
    SS3[0][47] = 4'h0;
    SS3[1][47] = 4'h0;
    SS3[2][47] = 4'h0;
    SS3[3][47] = 4'h0;
    SS3[4][47] = 4'h0;
    SS3[5][47] = 4'h0;
    SS3[6][47] = 4'h0;
    SS3[7][47] = 4'h0;
    SS3[8][47] = 4'h0;
    SS3[9][47] = 4'h0;
    SS3[10][47] = 4'h0;
    SS3[11][47] = 4'h0;
    SS3[12][47] = 4'h0;
    SS3[13][47] = 4'h0;
    SS3[14][47] = 4'h0;
    SS3[15][47] = 4'h0;
    SS3[16][47] = 4'h0;
    SS3[17][47] = 4'h0;
    SS3[18][47] = 4'h0;
    SS3[19][47] = 4'h0;
    SS3[20][47] = 4'h0;
    SS3[21][47] = 4'h0;
    SS3[22][47] = 4'h0;
    SS3[23][47] = 4'h0;
    SS3[24][47] = 4'hD;
    SS3[25][47] = 4'hD;
    SS3[26][47] = 4'hD;
    SS3[27][47] = 4'h0;
    SS3[28][47] = 4'h0;
    SS3[29][47] = 4'h0;
    SS3[30][47] = 4'h0;
    SS3[31][47] = 4'h0;
    SS3[32][47] = 4'h0;
    SS3[33][47] = 4'h0;
    SS3[34][47] = 4'h0;
    SS3[35][47] = 4'h0;
    SS3[36][47] = 4'h0;
    SS3[37][47] = 4'h0;
    SS3[38][47] = 4'h0;
    SS3[39][47] = 4'h0;
    SS3[40][47] = 4'h0;
    SS3[41][47] = 4'h0;
    SS3[42][47] = 4'h0;
    SS3[43][47] = 4'h0;
    SS3[44][47] = 4'h0;
    SS3[45][47] = 4'h0;
    SS3[46][47] = 4'h0;
    SS3[47][47] = 4'h0;
 
//SS 4
    SS4[0][0] = 4'h0;
    SS4[1][0] = 4'h0;
    SS4[2][0] = 4'h0;
    SS4[3][0] = 4'h0;
    SS4[4][0] = 4'h0;
    SS4[5][0] = 4'h0;
    SS4[6][0] = 4'h0;
    SS4[7][0] = 4'h0;
    SS4[8][0] = 4'h0;
    SS4[9][0] = 4'h0;
    SS4[10][0] = 4'h0;
    SS4[11][0] = 4'h0;
    SS4[12][0] = 4'h0;
    SS4[13][0] = 4'h0;
    SS4[14][0] = 4'h0;
    SS4[15][0] = 4'hD;
    SS4[16][0] = 4'hD;
    SS4[17][0] = 4'hD;
    SS4[18][0] = 4'h0;
    SS4[19][0] = 4'h0;
    SS4[20][0] = 4'h0;
    SS4[21][0] = 4'h0;
    SS4[22][0] = 4'h0;
    SS4[23][0] = 4'h0;
    SS4[24][0] = 4'h0;
    SS4[25][0] = 4'h0;
    SS4[26][0] = 4'h0;
    SS4[27][0] = 4'h0;
    SS4[28][0] = 4'h0;
    SS4[29][0] = 4'h0;
    SS4[30][0] = 4'h0;
    SS4[31][0] = 4'h0;
    SS4[32][0] = 4'h0;
    SS4[33][0] = 4'h0;
    SS4[34][0] = 4'h0;
    SS4[35][0] = 4'h0;
    SS4[36][0] = 4'h0;
    SS4[37][0] = 4'h0;
    SS4[38][0] = 4'h0;
    SS4[39][0] = 4'h0;
    SS4[40][0] = 4'h0;
    SS4[41][0] = 4'h0;
    SS4[42][0] = 4'h0;
    SS4[43][0] = 4'h0;
    SS4[44][0] = 4'h0;
    SS4[45][0] = 4'h0;
    SS4[46][0] = 4'h0;
    SS4[47][0] = 4'h0;
    SS4[0][1] = 4'h0;
    SS4[1][1] = 4'h0;
    SS4[2][1] = 4'h0;
    SS4[3][1] = 4'h0;
    SS4[4][1] = 4'h0;
    SS4[5][1] = 4'h0;
    SS4[6][1] = 4'h0;
    SS4[7][1] = 4'h0;
    SS4[8][1] = 4'h0;
    SS4[9][1] = 4'h0;
    SS4[10][1] = 4'h0;
    SS4[11][1] = 4'h0;
    SS4[12][1] = 4'h0;
    SS4[13][1] = 4'h0;
    SS4[14][1] = 4'h0;
    SS4[15][1] = 4'hD;
    SS4[16][1] = 4'hD;
    SS4[17][1] = 4'hD;
    SS4[18][1] = 4'h0;
    SS4[19][1] = 4'h0;
    SS4[20][1] = 4'h0;
    SS4[21][1] = 4'h0;
    SS4[22][1] = 4'h0;
    SS4[23][1] = 4'h0;
    SS4[24][1] = 4'h0;
    SS4[25][1] = 4'h0;
    SS4[26][1] = 4'h0;
    SS4[27][1] = 4'h0;
    SS4[28][1] = 4'h0;
    SS4[29][1] = 4'h0;
    SS4[30][1] = 4'h0;
    SS4[31][1] = 4'h0;
    SS4[32][1] = 4'h0;
    SS4[33][1] = 4'h0;
    SS4[34][1] = 4'h0;
    SS4[35][1] = 4'h0;
    SS4[36][1] = 4'h0;
    SS4[37][1] = 4'h0;
    SS4[38][1] = 4'h0;
    SS4[39][1] = 4'h0;
    SS4[40][1] = 4'h0;
    SS4[41][1] = 4'h0;
    SS4[42][1] = 4'h0;
    SS4[43][1] = 4'h0;
    SS4[44][1] = 4'h0;
    SS4[45][1] = 4'h0;
    SS4[46][1] = 4'h0;
    SS4[47][1] = 4'h0;
    SS4[0][2] = 4'h0;
    SS4[1][2] = 4'h0;
    SS4[2][2] = 4'h0;
    SS4[3][2] = 4'h0;
    SS4[4][2] = 4'h0;
    SS4[5][2] = 4'h0;
    SS4[6][2] = 4'h0;
    SS4[7][2] = 4'h0;
    SS4[8][2] = 4'h0;
    SS4[9][2] = 4'h0;
    SS4[10][2] = 4'h0;
    SS4[11][2] = 4'h0;
    SS4[12][2] = 4'h0;
    SS4[13][2] = 4'h0;
    SS4[14][2] = 4'h0;
    SS4[15][2] = 4'hD;
    SS4[16][2] = 4'hD;
    SS4[17][2] = 4'hD;
    SS4[18][2] = 4'h0;
    SS4[19][2] = 4'h0;
    SS4[20][2] = 4'h0;
    SS4[21][2] = 4'h0;
    SS4[22][2] = 4'h0;
    SS4[23][2] = 4'h0;
    SS4[24][2] = 4'h0;
    SS4[25][2] = 4'h0;
    SS4[26][2] = 4'h0;
    SS4[27][2] = 4'h0;
    SS4[28][2] = 4'h0;
    SS4[29][2] = 4'h0;
    SS4[30][2] = 4'h0;
    SS4[31][2] = 4'h0;
    SS4[32][2] = 4'h0;
    SS4[33][2] = 4'h0;
    SS4[34][2] = 4'h0;
    SS4[35][2] = 4'h0;
    SS4[36][2] = 4'h0;
    SS4[37][2] = 4'h0;
    SS4[38][2] = 4'h0;
    SS4[39][2] = 4'h0;
    SS4[40][2] = 4'h0;
    SS4[41][2] = 4'h0;
    SS4[42][2] = 4'h0;
    SS4[43][2] = 4'h0;
    SS4[44][2] = 4'h0;
    SS4[45][2] = 4'h0;
    SS4[46][2] = 4'h0;
    SS4[47][2] = 4'h0;
    SS4[0][3] = 4'h0;
    SS4[1][3] = 4'h0;
    SS4[2][3] = 4'h0;
    SS4[3][3] = 4'h0;
    SS4[4][3] = 4'h0;
    SS4[5][3] = 4'h0;
    SS4[6][3] = 4'h0;
    SS4[7][3] = 4'h0;
    SS4[8][3] = 4'h0;
    SS4[9][3] = 4'h0;
    SS4[10][3] = 4'h0;
    SS4[11][3] = 4'h0;
    SS4[12][3] = 4'h0;
    SS4[13][3] = 4'h0;
    SS4[14][3] = 4'h0;
    SS4[15][3] = 4'hD;
    SS4[16][3] = 4'hD;
    SS4[17][3] = 4'hD;
    SS4[18][3] = 4'hD;
    SS4[19][3] = 4'hD;
    SS4[20][3] = 4'hD;
    SS4[21][3] = 4'h0;
    SS4[22][3] = 4'h0;
    SS4[23][3] = 4'h0;
    SS4[24][3] = 4'h0;
    SS4[25][3] = 4'h0;
    SS4[26][3] = 4'h0;
    SS4[27][3] = 4'h0;
    SS4[28][3] = 4'h0;
    SS4[29][3] = 4'h0;
    SS4[30][3] = 4'h0;
    SS4[31][3] = 4'h0;
    SS4[32][3] = 4'h0;
    SS4[33][3] = 4'h0;
    SS4[34][3] = 4'h0;
    SS4[35][3] = 4'h0;
    SS4[36][3] = 4'h0;
    SS4[37][3] = 4'h0;
    SS4[38][3] = 4'h0;
    SS4[39][3] = 4'h0;
    SS4[40][3] = 4'h0;
    SS4[41][3] = 4'h0;
    SS4[42][3] = 4'h0;
    SS4[43][3] = 4'h0;
    SS4[44][3] = 4'h0;
    SS4[45][3] = 4'h0;
    SS4[46][3] = 4'h0;
    SS4[47][3] = 4'h0;
    SS4[0][4] = 4'h0;
    SS4[1][4] = 4'h0;
    SS4[2][4] = 4'h0;
    SS4[3][4] = 4'h0;
    SS4[4][4] = 4'h0;
    SS4[5][4] = 4'h0;
    SS4[6][4] = 4'h0;
    SS4[7][4] = 4'h0;
    SS4[8][4] = 4'h0;
    SS4[9][4] = 4'h0;
    SS4[10][4] = 4'h0;
    SS4[11][4] = 4'h0;
    SS4[12][4] = 4'h0;
    SS4[13][4] = 4'h0;
    SS4[14][4] = 4'h0;
    SS4[15][4] = 4'hD;
    SS4[16][4] = 4'hD;
    SS4[17][4] = 4'hD;
    SS4[18][4] = 4'hD;
    SS4[19][4] = 4'hD;
    SS4[20][4] = 4'hD;
    SS4[21][4] = 4'h0;
    SS4[22][4] = 4'h0;
    SS4[23][4] = 4'h0;
    SS4[24][4] = 4'h0;
    SS4[25][4] = 4'h0;
    SS4[26][4] = 4'h0;
    SS4[27][4] = 4'h0;
    SS4[28][4] = 4'h0;
    SS4[29][4] = 4'h0;
    SS4[30][4] = 4'h0;
    SS4[31][4] = 4'h0;
    SS4[32][4] = 4'h0;
    SS4[33][4] = 4'h0;
    SS4[34][4] = 4'h0;
    SS4[35][4] = 4'h0;
    SS4[36][4] = 4'h0;
    SS4[37][4] = 4'h0;
    SS4[38][4] = 4'h0;
    SS4[39][4] = 4'h0;
    SS4[40][4] = 4'h0;
    SS4[41][4] = 4'h0;
    SS4[42][4] = 4'h0;
    SS4[43][4] = 4'h0;
    SS4[44][4] = 4'h0;
    SS4[45][4] = 4'h0;
    SS4[46][4] = 4'h0;
    SS4[47][4] = 4'h0;
    SS4[0][5] = 4'h0;
    SS4[1][5] = 4'h0;
    SS4[2][5] = 4'h0;
    SS4[3][5] = 4'h0;
    SS4[4][5] = 4'h0;
    SS4[5][5] = 4'h0;
    SS4[6][5] = 4'h0;
    SS4[7][5] = 4'h0;
    SS4[8][5] = 4'h0;
    SS4[9][5] = 4'h0;
    SS4[10][5] = 4'h0;
    SS4[11][5] = 4'h0;
    SS4[12][5] = 4'h0;
    SS4[13][5] = 4'h0;
    SS4[14][5] = 4'h0;
    SS4[15][5] = 4'hD;
    SS4[16][5] = 4'hD;
    SS4[17][5] = 4'hD;
    SS4[18][5] = 4'hD;
    SS4[19][5] = 4'hD;
    SS4[20][5] = 4'hD;
    SS4[21][5] = 4'h0;
    SS4[22][5] = 4'h0;
    SS4[23][5] = 4'h0;
    SS4[24][5] = 4'h0;
    SS4[25][5] = 4'h0;
    SS4[26][5] = 4'h0;
    SS4[27][5] = 4'h0;
    SS4[28][5] = 4'h0;
    SS4[29][5] = 4'h0;
    SS4[30][5] = 4'h0;
    SS4[31][5] = 4'h0;
    SS4[32][5] = 4'h0;
    SS4[33][5] = 4'h0;
    SS4[34][5] = 4'h0;
    SS4[35][5] = 4'h0;
    SS4[36][5] = 4'h0;
    SS4[37][5] = 4'h0;
    SS4[38][5] = 4'h0;
    SS4[39][5] = 4'h0;
    SS4[40][5] = 4'h0;
    SS4[41][5] = 4'h0;
    SS4[42][5] = 4'h0;
    SS4[43][5] = 4'h0;
    SS4[44][5] = 4'h0;
    SS4[45][5] = 4'h0;
    SS4[46][5] = 4'h0;
    SS4[47][5] = 4'h0;
    SS4[0][6] = 4'h0;
    SS4[1][6] = 4'h0;
    SS4[2][6] = 4'h0;
    SS4[3][6] = 4'h0;
    SS4[4][6] = 4'h0;
    SS4[5][6] = 4'h0;
    SS4[6][6] = 4'h0;
    SS4[7][6] = 4'h0;
    SS4[8][6] = 4'h0;
    SS4[9][6] = 4'h0;
    SS4[10][6] = 4'h0;
    SS4[11][6] = 4'h0;
    SS4[12][6] = 4'h0;
    SS4[13][6] = 4'h0;
    SS4[14][6] = 4'h0;
    SS4[15][6] = 4'hE;
    SS4[16][6] = 4'hE;
    SS4[17][6] = 4'hE;
    SS4[18][6] = 4'hD;
    SS4[19][6] = 4'hD;
    SS4[20][6] = 4'hD;
    SS4[21][6] = 4'h3;
    SS4[22][6] = 4'h3;
    SS4[23][6] = 4'h3;
    SS4[24][6] = 4'h0;
    SS4[25][6] = 4'h0;
    SS4[26][6] = 4'h0;
    SS4[27][6] = 4'h0;
    SS4[28][6] = 4'h0;
    SS4[29][6] = 4'h0;
    SS4[30][6] = 4'h0;
    SS4[31][6] = 4'h0;
    SS4[32][6] = 4'h0;
    SS4[33][6] = 4'h0;
    SS4[34][6] = 4'h0;
    SS4[35][6] = 4'h0;
    SS4[36][6] = 4'h0;
    SS4[37][6] = 4'h0;
    SS4[38][6] = 4'h0;
    SS4[39][6] = 4'h0;
    SS4[40][6] = 4'h0;
    SS4[41][6] = 4'h0;
    SS4[42][6] = 4'h0;
    SS4[43][6] = 4'h0;
    SS4[44][6] = 4'h0;
    SS4[45][6] = 4'h0;
    SS4[46][6] = 4'h0;
    SS4[47][6] = 4'h0;
    SS4[0][7] = 4'h0;
    SS4[1][7] = 4'h0;
    SS4[2][7] = 4'h0;
    SS4[3][7] = 4'h0;
    SS4[4][7] = 4'h0;
    SS4[5][7] = 4'h0;
    SS4[6][7] = 4'h0;
    SS4[7][7] = 4'h0;
    SS4[8][7] = 4'h0;
    SS4[9][7] = 4'h0;
    SS4[10][7] = 4'h0;
    SS4[11][7] = 4'h0;
    SS4[12][7] = 4'h0;
    SS4[13][7] = 4'h0;
    SS4[14][7] = 4'h0;
    SS4[15][7] = 4'hE;
    SS4[16][7] = 4'hE;
    SS4[17][7] = 4'hE;
    SS4[18][7] = 4'hD;
    SS4[19][7] = 4'hD;
    SS4[20][7] = 4'hD;
    SS4[21][7] = 4'h3;
    SS4[22][7] = 4'h3;
    SS4[23][7] = 4'h3;
    SS4[24][7] = 4'h0;
    SS4[25][7] = 4'h0;
    SS4[26][7] = 4'h0;
    SS4[27][7] = 4'h0;
    SS4[28][7] = 4'h0;
    SS4[29][7] = 4'h0;
    SS4[30][7] = 4'h0;
    SS4[31][7] = 4'h0;
    SS4[32][7] = 4'h0;
    SS4[33][7] = 4'h0;
    SS4[34][7] = 4'h0;
    SS4[35][7] = 4'h0;
    SS4[36][7] = 4'h0;
    SS4[37][7] = 4'h0;
    SS4[38][7] = 4'h0;
    SS4[39][7] = 4'h0;
    SS4[40][7] = 4'h0;
    SS4[41][7] = 4'h0;
    SS4[42][7] = 4'h0;
    SS4[43][7] = 4'h0;
    SS4[44][7] = 4'h0;
    SS4[45][7] = 4'h0;
    SS4[46][7] = 4'h0;
    SS4[47][7] = 4'h0;
    SS4[0][8] = 4'h0;
    SS4[1][8] = 4'h0;
    SS4[2][8] = 4'h0;
    SS4[3][8] = 4'h0;
    SS4[4][8] = 4'h0;
    SS4[5][8] = 4'h0;
    SS4[6][8] = 4'h0;
    SS4[7][8] = 4'h0;
    SS4[8][8] = 4'h0;
    SS4[9][8] = 4'h0;
    SS4[10][8] = 4'h0;
    SS4[11][8] = 4'h0;
    SS4[12][8] = 4'h0;
    SS4[13][8] = 4'h0;
    SS4[14][8] = 4'h0;
    SS4[15][8] = 4'hE;
    SS4[16][8] = 4'hE;
    SS4[17][8] = 4'hE;
    SS4[18][8] = 4'hD;
    SS4[19][8] = 4'hD;
    SS4[20][8] = 4'hD;
    SS4[21][8] = 4'h3;
    SS4[22][8] = 4'h3;
    SS4[23][8] = 4'h3;
    SS4[24][8] = 4'h0;
    SS4[25][8] = 4'h0;
    SS4[26][8] = 4'h0;
    SS4[27][8] = 4'h0;
    SS4[28][8] = 4'h0;
    SS4[29][8] = 4'h0;
    SS4[30][8] = 4'h0;
    SS4[31][8] = 4'h0;
    SS4[32][8] = 4'h0;
    SS4[33][8] = 4'h0;
    SS4[34][8] = 4'h0;
    SS4[35][8] = 4'h0;
    SS4[36][8] = 4'h0;
    SS4[37][8] = 4'h0;
    SS4[38][8] = 4'h0;
    SS4[39][8] = 4'h0;
    SS4[40][8] = 4'h0;
    SS4[41][8] = 4'h0;
    SS4[42][8] = 4'h0;
    SS4[43][8] = 4'h0;
    SS4[44][8] = 4'h0;
    SS4[45][8] = 4'h0;
    SS4[46][8] = 4'h0;
    SS4[47][8] = 4'h0;
    SS4[0][9] = 4'hD;
    SS4[1][9] = 4'hD;
    SS4[2][9] = 4'hD;
    SS4[3][9] = 4'hC;
    SS4[4][9] = 4'hC;
    SS4[5][9] = 4'hC;
    SS4[6][9] = 4'hC;
    SS4[7][9] = 4'hC;
    SS4[8][9] = 4'hC;
    SS4[9][9] = 4'h0;
    SS4[10][9] = 4'h0;
    SS4[11][9] = 4'h0;
    SS4[12][9] = 4'h0;
    SS4[13][9] = 4'h0;
    SS4[14][9] = 4'h0;
    SS4[15][9] = 4'hE;
    SS4[16][9] = 4'hE;
    SS4[17][9] = 4'hE;
    SS4[18][9] = 4'hE;
    SS4[19][9] = 4'hE;
    SS4[20][9] = 4'hE;
    SS4[21][9] = 4'hD;
    SS4[22][9] = 4'hD;
    SS4[23][9] = 4'hD;
    SS4[24][9] = 4'h0;
    SS4[25][9] = 4'h0;
    SS4[26][9] = 4'h0;
    SS4[27][9] = 4'h0;
    SS4[28][9] = 4'h0;
    SS4[29][9] = 4'h0;
    SS4[30][9] = 4'h0;
    SS4[31][9] = 4'h0;
    SS4[32][9] = 4'h0;
    SS4[33][9] = 4'h0;
    SS4[34][9] = 4'h0;
    SS4[35][9] = 4'h0;
    SS4[36][9] = 4'h0;
    SS4[37][9] = 4'h0;
    SS4[38][9] = 4'h0;
    SS4[39][9] = 4'h0;
    SS4[40][9] = 4'h0;
    SS4[41][9] = 4'h0;
    SS4[42][9] = 4'h0;
    SS4[43][9] = 4'h0;
    SS4[44][9] = 4'h0;
    SS4[45][9] = 4'h0;
    SS4[46][9] = 4'h0;
    SS4[47][9] = 4'h0;
    SS4[0][10] = 4'hD;
    SS4[1][10] = 4'hD;
    SS4[2][10] = 4'hD;
    SS4[3][10] = 4'hC;
    SS4[4][10] = 4'hC;
    SS4[5][10] = 4'hC;
    SS4[6][10] = 4'hC;
    SS4[7][10] = 4'hC;
    SS4[8][10] = 4'hC;
    SS4[9][10] = 4'h0;
    SS4[10][10] = 4'h0;
    SS4[11][10] = 4'h0;
    SS4[12][10] = 4'h0;
    SS4[13][10] = 4'h0;
    SS4[14][10] = 4'h0;
    SS4[15][10] = 4'hE;
    SS4[16][10] = 4'hE;
    SS4[17][10] = 4'hE;
    SS4[18][10] = 4'hE;
    SS4[19][10] = 4'hE;
    SS4[20][10] = 4'hE;
    SS4[21][10] = 4'hD;
    SS4[22][10] = 4'hD;
    SS4[23][10] = 4'hD;
    SS4[24][10] = 4'h0;
    SS4[25][10] = 4'h0;
    SS4[26][10] = 4'h0;
    SS4[27][10] = 4'h0;
    SS4[28][10] = 4'h0;
    SS4[29][10] = 4'h0;
    SS4[30][10] = 4'h0;
    SS4[31][10] = 4'h0;
    SS4[32][10] = 4'h0;
    SS4[33][10] = 4'h0;
    SS4[34][10] = 4'h0;
    SS4[35][10] = 4'h0;
    SS4[36][10] = 4'h0;
    SS4[37][10] = 4'h0;
    SS4[38][10] = 4'h0;
    SS4[39][10] = 4'h0;
    SS4[40][10] = 4'h0;
    SS4[41][10] = 4'h0;
    SS4[42][10] = 4'h0;
    SS4[43][10] = 4'h0;
    SS4[44][10] = 4'h0;
    SS4[45][10] = 4'h0;
    SS4[46][10] = 4'h0;
    SS4[47][10] = 4'h0;
    SS4[0][11] = 4'hD;
    SS4[1][11] = 4'hD;
    SS4[2][11] = 4'hD;
    SS4[3][11] = 4'hC;
    SS4[4][11] = 4'hC;
    SS4[5][11] = 4'hC;
    SS4[6][11] = 4'hC;
    SS4[7][11] = 4'hC;
    SS4[8][11] = 4'hC;
    SS4[9][11] = 4'h0;
    SS4[10][11] = 4'h0;
    SS4[11][11] = 4'h0;
    SS4[12][11] = 4'h0;
    SS4[13][11] = 4'h0;
    SS4[14][11] = 4'h0;
    SS4[15][11] = 4'hE;
    SS4[16][11] = 4'hE;
    SS4[17][11] = 4'hE;
    SS4[18][11] = 4'hE;
    SS4[19][11] = 4'hE;
    SS4[20][11] = 4'hE;
    SS4[21][11] = 4'hD;
    SS4[22][11] = 4'hD;
    SS4[23][11] = 4'hD;
    SS4[24][11] = 4'h0;
    SS4[25][11] = 4'h0;
    SS4[26][11] = 4'h0;
    SS4[27][11] = 4'h0;
    SS4[28][11] = 4'h0;
    SS4[29][11] = 4'h0;
    SS4[30][11] = 4'h0;
    SS4[31][11] = 4'h0;
    SS4[32][11] = 4'h0;
    SS4[33][11] = 4'h0;
    SS4[34][11] = 4'h0;
    SS4[35][11] = 4'h0;
    SS4[36][11] = 4'h0;
    SS4[37][11] = 4'h0;
    SS4[38][11] = 4'h0;
    SS4[39][11] = 4'h0;
    SS4[40][11] = 4'h0;
    SS4[41][11] = 4'h0;
    SS4[42][11] = 4'h0;
    SS4[43][11] = 4'h0;
    SS4[44][11] = 4'h0;
    SS4[45][11] = 4'h0;
    SS4[46][11] = 4'h0;
    SS4[47][11] = 4'h0;
    SS4[0][12] = 4'h0;
    SS4[1][12] = 4'h0;
    SS4[2][12] = 4'h0;
    SS4[3][12] = 4'hD;
    SS4[4][12] = 4'hD;
    SS4[5][12] = 4'hD;
    SS4[6][12] = 4'hC;
    SS4[7][12] = 4'hC;
    SS4[8][12] = 4'hC;
    SS4[9][12] = 4'hC;
    SS4[10][12] = 4'hC;
    SS4[11][12] = 4'hC;
    SS4[12][12] = 4'hC;
    SS4[13][12] = 4'hC;
    SS4[14][12] = 4'hC;
    SS4[15][12] = 4'hC;
    SS4[16][12] = 4'hC;
    SS4[17][12] = 4'hC;
    SS4[18][12] = 4'hE;
    SS4[19][12] = 4'hE;
    SS4[20][12] = 4'hE;
    SS4[21][12] = 4'hD;
    SS4[22][12] = 4'hD;
    SS4[23][12] = 4'hD;
    SS4[24][12] = 4'hD;
    SS4[25][12] = 4'hD;
    SS4[26][12] = 4'hD;
    SS4[27][12] = 4'h3;
    SS4[28][12] = 4'h3;
    SS4[29][12] = 4'h3;
    SS4[30][12] = 4'h0;
    SS4[31][12] = 4'h0;
    SS4[32][12] = 4'h0;
    SS4[33][12] = 4'h0;
    SS4[34][12] = 4'h0;
    SS4[35][12] = 4'h0;
    SS4[36][12] = 4'h0;
    SS4[37][12] = 4'h0;
    SS4[38][12] = 4'h0;
    SS4[39][12] = 4'h0;
    SS4[40][12] = 4'h0;
    SS4[41][12] = 4'h0;
    SS4[42][12] = 4'h0;
    SS4[43][12] = 4'h0;
    SS4[44][12] = 4'h0;
    SS4[45][12] = 4'h0;
    SS4[46][12] = 4'h0;
    SS4[47][12] = 4'h0;
    SS4[0][13] = 4'h0;
    SS4[1][13] = 4'h0;
    SS4[2][13] = 4'h0;
    SS4[3][13] = 4'hD;
    SS4[4][13] = 4'hD;
    SS4[5][13] = 4'hD;
    SS4[6][13] = 4'hC;
    SS4[7][13] = 4'hC;
    SS4[8][13] = 4'hC;
    SS4[9][13] = 4'hC;
    SS4[10][13] = 4'hC;
    SS4[11][13] = 4'hC;
    SS4[12][13] = 4'hC;
    SS4[13][13] = 4'hC;
    SS4[14][13] = 4'hC;
    SS4[15][13] = 4'hC;
    SS4[16][13] = 4'hC;
    SS4[17][13] = 4'hC;
    SS4[18][13] = 4'hE;
    SS4[19][13] = 4'hE;
    SS4[20][13] = 4'hE;
    SS4[21][13] = 4'hD;
    SS4[22][13] = 4'hD;
    SS4[23][13] = 4'hD;
    SS4[24][13] = 4'hD;
    SS4[25][13] = 4'hD;
    SS4[26][13] = 4'hD;
    SS4[27][13] = 4'h3;
    SS4[28][13] = 4'h3;
    SS4[29][13] = 4'h3;
    SS4[30][13] = 4'h0;
    SS4[31][13] = 4'h0;
    SS4[32][13] = 4'h0;
    SS4[33][13] = 4'h0;
    SS4[34][13] = 4'h0;
    SS4[35][13] = 4'h0;
    SS4[36][13] = 4'h0;
    SS4[37][13] = 4'h0;
    SS4[38][13] = 4'h0;
    SS4[39][13] = 4'h0;
    SS4[40][13] = 4'h0;
    SS4[41][13] = 4'h0;
    SS4[42][13] = 4'h0;
    SS4[43][13] = 4'h0;
    SS4[44][13] = 4'h0;
    SS4[45][13] = 4'h0;
    SS4[46][13] = 4'h0;
    SS4[47][13] = 4'h0;
    SS4[0][14] = 4'h0;
    SS4[1][14] = 4'h0;
    SS4[2][14] = 4'h0;
    SS4[3][14] = 4'hD;
    SS4[4][14] = 4'hD;
    SS4[5][14] = 4'hD;
    SS4[6][14] = 4'hC;
    SS4[7][14] = 4'hC;
    SS4[8][14] = 4'hC;
    SS4[9][14] = 4'hC;
    SS4[10][14] = 4'hC;
    SS4[11][14] = 4'hC;
    SS4[12][14] = 4'hC;
    SS4[13][14] = 4'hC;
    SS4[14][14] = 4'hC;
    SS4[15][14] = 4'hC;
    SS4[16][14] = 4'hC;
    SS4[17][14] = 4'hC;
    SS4[18][14] = 4'hE;
    SS4[19][14] = 4'hE;
    SS4[20][14] = 4'hE;
    SS4[21][14] = 4'hD;
    SS4[22][14] = 4'hD;
    SS4[23][14] = 4'hD;
    SS4[24][14] = 4'hD;
    SS4[25][14] = 4'hD;
    SS4[26][14] = 4'hD;
    SS4[27][14] = 4'h3;
    SS4[28][14] = 4'h3;
    SS4[29][14] = 4'h3;
    SS4[30][14] = 4'h0;
    SS4[31][14] = 4'h0;
    SS4[32][14] = 4'h0;
    SS4[33][14] = 4'h0;
    SS4[34][14] = 4'h0;
    SS4[35][14] = 4'h0;
    SS4[36][14] = 4'h0;
    SS4[37][14] = 4'h0;
    SS4[38][14] = 4'h0;
    SS4[39][14] = 4'h0;
    SS4[40][14] = 4'h0;
    SS4[41][14] = 4'h0;
    SS4[42][14] = 4'h0;
    SS4[43][14] = 4'h0;
    SS4[44][14] = 4'h0;
    SS4[45][14] = 4'h0;
    SS4[46][14] = 4'h0;
    SS4[47][14] = 4'h0;
    SS4[0][15] = 4'h0;
    SS4[1][15] = 4'h0;
    SS4[2][15] = 4'h0;
    SS4[3][15] = 4'h0;
    SS4[4][15] = 4'h0;
    SS4[5][15] = 4'h0;
    SS4[6][15] = 4'hE;
    SS4[7][15] = 4'hE;
    SS4[8][15] = 4'hE;
    SS4[9][15] = 4'hD;
    SS4[10][15] = 4'hD;
    SS4[11][15] = 4'hD;
    SS4[12][15] = 4'hC;
    SS4[13][15] = 4'hC;
    SS4[14][15] = 4'hC;
    SS4[15][15] = 4'hC;
    SS4[16][15] = 4'hC;
    SS4[17][15] = 4'hC;
    SS4[18][15] = 4'hC;
    SS4[19][15] = 4'hC;
    SS4[20][15] = 4'hC;
    SS4[21][15] = 4'hE;
    SS4[22][15] = 4'hE;
    SS4[23][15] = 4'hE;
    SS4[24][15] = 4'hD;
    SS4[25][15] = 4'hD;
    SS4[26][15] = 4'hD;
    SS4[27][15] = 4'hD;
    SS4[28][15] = 4'hD;
    SS4[29][15] = 4'hD;
    SS4[30][15] = 4'h0;
    SS4[31][15] = 4'h0;
    SS4[32][15] = 4'h0;
    SS4[33][15] = 4'h0;
    SS4[34][15] = 4'h0;
    SS4[35][15] = 4'h0;
    SS4[36][15] = 4'h0;
    SS4[37][15] = 4'h0;
    SS4[38][15] = 4'h0;
    SS4[39][15] = 4'h0;
    SS4[40][15] = 4'h0;
    SS4[41][15] = 4'h0;
    SS4[42][15] = 4'h0;
    SS4[43][15] = 4'h0;
    SS4[44][15] = 4'h0;
    SS4[45][15] = 4'h0;
    SS4[46][15] = 4'h0;
    SS4[47][15] = 4'h0;
    SS4[0][16] = 4'h0;
    SS4[1][16] = 4'h0;
    SS4[2][16] = 4'h0;
    SS4[3][16] = 4'h0;
    SS4[4][16] = 4'h0;
    SS4[5][16] = 4'h0;
    SS4[6][16] = 4'hE;
    SS4[7][16] = 4'hE;
    SS4[8][16] = 4'hE;
    SS4[9][16] = 4'hD;
    SS4[10][16] = 4'hD;
    SS4[11][16] = 4'hD;
    SS4[12][16] = 4'hC;
    SS4[13][16] = 4'hC;
    SS4[14][16] = 4'hC;
    SS4[15][16] = 4'hC;
    SS4[16][16] = 4'hC;
    SS4[17][16] = 4'hC;
    SS4[18][16] = 4'hC;
    SS4[19][16] = 4'hC;
    SS4[20][16] = 4'hC;
    SS4[21][16] = 4'hE;
    SS4[22][16] = 4'hE;
    SS4[23][16] = 4'hE;
    SS4[24][16] = 4'hD;
    SS4[25][16] = 4'hD;
    SS4[26][16] = 4'hD;
    SS4[27][16] = 4'hD;
    SS4[28][16] = 4'hD;
    SS4[29][16] = 4'hD;
    SS4[30][16] = 4'h0;
    SS4[31][16] = 4'h0;
    SS4[32][16] = 4'h0;
    SS4[33][16] = 4'h0;
    SS4[34][16] = 4'h0;
    SS4[35][16] = 4'h0;
    SS4[36][16] = 4'h0;
    SS4[37][16] = 4'h0;
    SS4[38][16] = 4'h0;
    SS4[39][16] = 4'h0;
    SS4[40][16] = 4'h0;
    SS4[41][16] = 4'h0;
    SS4[42][16] = 4'h0;
    SS4[43][16] = 4'h0;
    SS4[44][16] = 4'h0;
    SS4[45][16] = 4'h0;
    SS4[46][16] = 4'h0;
    SS4[47][16] = 4'h0;
    SS4[0][17] = 4'h0;
    SS4[1][17] = 4'h0;
    SS4[2][17] = 4'h0;
    SS4[3][17] = 4'h0;
    SS4[4][17] = 4'h0;
    SS4[5][17] = 4'h0;
    SS4[6][17] = 4'hE;
    SS4[7][17] = 4'hE;
    SS4[8][17] = 4'hE;
    SS4[9][17] = 4'hD;
    SS4[10][17] = 4'hD;
    SS4[11][17] = 4'hD;
    SS4[12][17] = 4'hC;
    SS4[13][17] = 4'hC;
    SS4[14][17] = 4'hC;
    SS4[15][17] = 4'hC;
    SS4[16][17] = 4'hC;
    SS4[17][17] = 4'hC;
    SS4[18][17] = 4'hC;
    SS4[19][17] = 4'hC;
    SS4[20][17] = 4'hC;
    SS4[21][17] = 4'hE;
    SS4[22][17] = 4'hE;
    SS4[23][17] = 4'hE;
    SS4[24][17] = 4'hD;
    SS4[25][17] = 4'hD;
    SS4[26][17] = 4'hD;
    SS4[27][17] = 4'hD;
    SS4[28][17] = 4'hD;
    SS4[29][17] = 4'hD;
    SS4[30][17] = 4'h0;
    SS4[31][17] = 4'h0;
    SS4[32][17] = 4'h0;
    SS4[33][17] = 4'h0;
    SS4[34][17] = 4'h0;
    SS4[35][17] = 4'h0;
    SS4[36][17] = 4'h0;
    SS4[37][17] = 4'h0;
    SS4[38][17] = 4'h0;
    SS4[39][17] = 4'h0;
    SS4[40][17] = 4'h0;
    SS4[41][17] = 4'h0;
    SS4[42][17] = 4'h0;
    SS4[43][17] = 4'h0;
    SS4[44][17] = 4'h0;
    SS4[45][17] = 4'h0;
    SS4[46][17] = 4'h0;
    SS4[47][17] = 4'h0;
    SS4[0][18] = 4'h0;
    SS4[1][18] = 4'h0;
    SS4[2][18] = 4'h0;
    SS4[3][18] = 4'h0;
    SS4[4][18] = 4'h0;
    SS4[5][18] = 4'h0;
    SS4[6][18] = 4'h0;
    SS4[7][18] = 4'h0;
    SS4[8][18] = 4'h0;
    SS4[9][18] = 4'hE;
    SS4[10][18] = 4'hE;
    SS4[11][18] = 4'hE;
    SS4[12][18] = 4'hD;
    SS4[13][18] = 4'hD;
    SS4[14][18] = 4'hD;
    SS4[15][18] = 4'hC;
    SS4[16][18] = 4'hC;
    SS4[17][18] = 4'hC;
    SS4[18][18] = 4'hC;
    SS4[19][18] = 4'hC;
    SS4[20][18] = 4'hC;
    SS4[21][18] = 4'hC;
    SS4[22][18] = 4'hC;
    SS4[23][18] = 4'hC;
    SS4[24][18] = 4'hC;
    SS4[25][18] = 4'hC;
    SS4[26][18] = 4'hC;
    SS4[27][18] = 4'hD;
    SS4[28][18] = 4'hD;
    SS4[29][18] = 4'hD;
    SS4[30][18] = 4'hC;
    SS4[31][18] = 4'hC;
    SS4[32][18] = 4'hC;
    SS4[33][18] = 4'hD;
    SS4[34][18] = 4'hD;
    SS4[35][18] = 4'hD;
    SS4[36][18] = 4'hD;
    SS4[37][18] = 4'hD;
    SS4[38][18] = 4'hD;
    SS4[39][18] = 4'hD;
    SS4[40][18] = 4'hD;
    SS4[41][18] = 4'hD;
    SS4[42][18] = 4'h0;
    SS4[43][18] = 4'h0;
    SS4[44][18] = 4'h0;
    SS4[45][18] = 4'h0;
    SS4[46][18] = 4'h0;
    SS4[47][18] = 4'h0;
    SS4[0][19] = 4'h0;
    SS4[1][19] = 4'h0;
    SS4[2][19] = 4'h0;
    SS4[3][19] = 4'h0;
    SS4[4][19] = 4'h0;
    SS4[5][19] = 4'h0;
    SS4[6][19] = 4'h0;
    SS4[7][19] = 4'h0;
    SS4[8][19] = 4'h0;
    SS4[9][19] = 4'hE;
    SS4[10][19] = 4'hE;
    SS4[11][19] = 4'hE;
    SS4[12][19] = 4'hD;
    SS4[13][19] = 4'hD;
    SS4[14][19] = 4'hD;
    SS4[15][19] = 4'hC;
    SS4[16][19] = 4'hC;
    SS4[17][19] = 4'hC;
    SS4[18][19] = 4'hC;
    SS4[19][19] = 4'hC;
    SS4[20][19] = 4'hC;
    SS4[21][19] = 4'hC;
    SS4[22][19] = 4'hC;
    SS4[23][19] = 4'hC;
    SS4[24][19] = 4'hC;
    SS4[25][19] = 4'hC;
    SS4[26][19] = 4'hC;
    SS4[27][19] = 4'hD;
    SS4[28][19] = 4'hD;
    SS4[29][19] = 4'hD;
    SS4[30][19] = 4'hC;
    SS4[31][19] = 4'hC;
    SS4[32][19] = 4'hC;
    SS4[33][19] = 4'hD;
    SS4[34][19] = 4'hD;
    SS4[35][19] = 4'hD;
    SS4[36][19] = 4'hD;
    SS4[37][19] = 4'hD;
    SS4[38][19] = 4'hD;
    SS4[39][19] = 4'hD;
    SS4[40][19] = 4'hD;
    SS4[41][19] = 4'hD;
    SS4[42][19] = 4'h0;
    SS4[43][19] = 4'h0;
    SS4[44][19] = 4'h0;
    SS4[45][19] = 4'h0;
    SS4[46][19] = 4'h0;
    SS4[47][19] = 4'h0;
    SS4[0][20] = 4'h0;
    SS4[1][20] = 4'h0;
    SS4[2][20] = 4'h0;
    SS4[3][20] = 4'h0;
    SS4[4][20] = 4'h0;
    SS4[5][20] = 4'h0;
    SS4[6][20] = 4'h0;
    SS4[7][20] = 4'h0;
    SS4[8][20] = 4'h0;
    SS4[9][20] = 4'hE;
    SS4[10][20] = 4'hE;
    SS4[11][20] = 4'hE;
    SS4[12][20] = 4'hD;
    SS4[13][20] = 4'hD;
    SS4[14][20] = 4'hD;
    SS4[15][20] = 4'hC;
    SS4[16][20] = 4'hC;
    SS4[17][20] = 4'hC;
    SS4[18][20] = 4'hC;
    SS4[19][20] = 4'hC;
    SS4[20][20] = 4'hC;
    SS4[21][20] = 4'hC;
    SS4[22][20] = 4'hC;
    SS4[23][20] = 4'hC;
    SS4[24][20] = 4'hC;
    SS4[25][20] = 4'hC;
    SS4[26][20] = 4'hC;
    SS4[27][20] = 4'hD;
    SS4[28][20] = 4'hD;
    SS4[29][20] = 4'hD;
    SS4[30][20] = 4'hC;
    SS4[31][20] = 4'hC;
    SS4[32][20] = 4'hC;
    SS4[33][20] = 4'hD;
    SS4[34][20] = 4'hD;
    SS4[35][20] = 4'hD;
    SS4[36][20] = 4'hD;
    SS4[37][20] = 4'hD;
    SS4[38][20] = 4'hD;
    SS4[39][20] = 4'hD;
    SS4[40][20] = 4'hD;
    SS4[41][20] = 4'hD;
    SS4[42][20] = 4'h0;
    SS4[43][20] = 4'h0;
    SS4[44][20] = 4'h0;
    SS4[45][20] = 4'h0;
    SS4[46][20] = 4'h0;
    SS4[47][20] = 4'h0;
    SS4[0][21] = 4'h0;
    SS4[1][21] = 4'h0;
    SS4[2][21] = 4'h0;
    SS4[3][21] = 4'h0;
    SS4[4][21] = 4'h0;
    SS4[5][21] = 4'h0;
    SS4[6][21] = 4'h0;
    SS4[7][21] = 4'h0;
    SS4[8][21] = 4'h0;
    SS4[9][21] = 4'h0;
    SS4[10][21] = 4'h0;
    SS4[11][21] = 4'h0;
    SS4[12][21] = 4'hE;
    SS4[13][21] = 4'hE;
    SS4[14][21] = 4'hE;
    SS4[15][21] = 4'hE;
    SS4[16][21] = 4'hE;
    SS4[17][21] = 4'hE;
    SS4[18][21] = 4'hD;
    SS4[19][21] = 4'hD;
    SS4[20][21] = 4'hD;
    SS4[21][21] = 4'hC;
    SS4[22][21] = 4'hC;
    SS4[23][21] = 4'hC;
    SS4[24][21] = 4'hD;
    SS4[25][21] = 4'hD;
    SS4[26][21] = 4'hD;
    SS4[27][21] = 4'hA;
    SS4[28][21] = 4'hA;
    SS4[29][21] = 4'hA;
    SS4[30][21] = 4'hC;
    SS4[31][21] = 4'hC;
    SS4[32][21] = 4'hC;
    SS4[33][21] = 4'hC;
    SS4[34][21] = 4'hC;
    SS4[35][21] = 4'hC;
    SS4[36][21] = 4'hC;
    SS4[37][21] = 4'hC;
    SS4[38][21] = 4'hC;
    SS4[39][21] = 4'hC;
    SS4[40][21] = 4'hC;
    SS4[41][21] = 4'hC;
    SS4[42][21] = 4'hC;
    SS4[43][21] = 4'hC;
    SS4[44][21] = 4'hC;
    SS4[45][21] = 4'hC;
    SS4[46][21] = 4'hC;
    SS4[47][21] = 4'hC;
    SS4[0][22] = 4'h0;
    SS4[1][22] = 4'h0;
    SS4[2][22] = 4'h0;
    SS4[3][22] = 4'h0;
    SS4[4][22] = 4'h0;
    SS4[5][22] = 4'h0;
    SS4[6][22] = 4'h0;
    SS4[7][22] = 4'h0;
    SS4[8][22] = 4'h0;
    SS4[9][22] = 4'h0;
    SS4[10][22] = 4'h0;
    SS4[11][22] = 4'h0;
    SS4[12][22] = 4'hE;
    SS4[13][22] = 4'hE;
    SS4[14][22] = 4'hE;
    SS4[15][22] = 4'hE;
    SS4[16][22] = 4'hE;
    SS4[17][22] = 4'hE;
    SS4[18][22] = 4'hD;
    SS4[19][22] = 4'hD;
    SS4[20][22] = 4'hD;
    SS4[21][22] = 4'hC;
    SS4[22][22] = 4'hC;
    SS4[23][22] = 4'hC;
    SS4[24][22] = 4'hD;
    SS4[25][22] = 4'hD;
    SS4[26][22] = 4'hD;
    SS4[27][22] = 4'hA;
    SS4[28][22] = 4'hA;
    SS4[29][22] = 4'hA;
    SS4[30][22] = 4'hC;
    SS4[31][22] = 4'hC;
    SS4[32][22] = 4'hC;
    SS4[33][22] = 4'hC;
    SS4[34][22] = 4'hC;
    SS4[35][22] = 4'hC;
    SS4[36][22] = 4'hC;
    SS4[37][22] = 4'hC;
    SS4[38][22] = 4'hC;
    SS4[39][22] = 4'hC;
    SS4[40][22] = 4'hC;
    SS4[41][22] = 4'hC;
    SS4[42][22] = 4'hC;
    SS4[43][22] = 4'hC;
    SS4[44][22] = 4'hC;
    SS4[45][22] = 4'hC;
    SS4[46][22] = 4'hC;
    SS4[47][22] = 4'hC;
    SS4[0][23] = 4'h0;
    SS4[1][23] = 4'h0;
    SS4[2][23] = 4'h0;
    SS4[3][23] = 4'h0;
    SS4[4][23] = 4'h0;
    SS4[5][23] = 4'h0;
    SS4[6][23] = 4'h0;
    SS4[7][23] = 4'h0;
    SS4[8][23] = 4'h0;
    SS4[9][23] = 4'h0;
    SS4[10][23] = 4'h0;
    SS4[11][23] = 4'h0;
    SS4[12][23] = 4'hE;
    SS4[13][23] = 4'hE;
    SS4[14][23] = 4'hE;
    SS4[15][23] = 4'hE;
    SS4[16][23] = 4'hE;
    SS4[17][23] = 4'hE;
    SS4[18][23] = 4'hD;
    SS4[19][23] = 4'hD;
    SS4[20][23] = 4'hD;
    SS4[21][23] = 4'hC;
    SS4[22][23] = 4'hC;
    SS4[23][23] = 4'hC;
    SS4[24][23] = 4'hD;
    SS4[25][23] = 4'hD;
    SS4[26][23] = 4'hD;
    SS4[27][23] = 4'hA;
    SS4[28][23] = 4'hA;
    SS4[29][23] = 4'hA;
    SS4[30][23] = 4'hC;
    SS4[31][23] = 4'hC;
    SS4[32][23] = 4'hC;
    SS4[33][23] = 4'hC;
    SS4[34][23] = 4'hC;
    SS4[35][23] = 4'hC;
    SS4[36][23] = 4'hC;
    SS4[37][23] = 4'hC;
    SS4[38][23] = 4'hC;
    SS4[39][23] = 4'hC;
    SS4[40][23] = 4'hC;
    SS4[41][23] = 4'hC;
    SS4[42][23] = 4'hC;
    SS4[43][23] = 4'hC;
    SS4[44][23] = 4'hC;
    SS4[45][23] = 4'hC;
    SS4[46][23] = 4'hC;
    SS4[47][23] = 4'hC;
    SS4[0][24] = 4'h0;
    SS4[1][24] = 4'h0;
    SS4[2][24] = 4'h0;
    SS4[3][24] = 4'h0;
    SS4[4][24] = 4'h0;
    SS4[5][24] = 4'h0;
    SS4[6][24] = 4'h0;
    SS4[7][24] = 4'h0;
    SS4[8][24] = 4'h0;
    SS4[9][24] = 4'h0;
    SS4[10][24] = 4'h0;
    SS4[11][24] = 4'h0;
    SS4[12][24] = 4'hE;
    SS4[13][24] = 4'hE;
    SS4[14][24] = 4'hE;
    SS4[15][24] = 4'hE;
    SS4[16][24] = 4'hE;
    SS4[17][24] = 4'hE;
    SS4[18][24] = 4'hD;
    SS4[19][24] = 4'hD;
    SS4[20][24] = 4'hD;
    SS4[21][24] = 4'hC;
    SS4[22][24] = 4'hC;
    SS4[23][24] = 4'hC;
    SS4[24][24] = 4'hD;
    SS4[25][24] = 4'hD;
    SS4[26][24] = 4'hD;
    SS4[27][24] = 4'hA;
    SS4[28][24] = 4'hA;
    SS4[29][24] = 4'hA;
    SS4[30][24] = 4'hC;
    SS4[31][24] = 4'hC;
    SS4[32][24] = 4'hC;
    SS4[33][24] = 4'hC;
    SS4[34][24] = 4'hC;
    SS4[35][24] = 4'hC;
    SS4[36][24] = 4'hC;
    SS4[37][24] = 4'hC;
    SS4[38][24] = 4'hC;
    SS4[39][24] = 4'hC;
    SS4[40][24] = 4'hC;
    SS4[41][24] = 4'hC;
    SS4[42][24] = 4'hC;
    SS4[43][24] = 4'hC;
    SS4[44][24] = 4'hC;
    SS4[45][24] = 4'hC;
    SS4[46][24] = 4'hC;
    SS4[47][24] = 4'hC;
    SS4[0][25] = 4'h0;
    SS4[1][25] = 4'h0;
    SS4[2][25] = 4'h0;
    SS4[3][25] = 4'h0;
    SS4[4][25] = 4'h0;
    SS4[5][25] = 4'h0;
    SS4[6][25] = 4'h0;
    SS4[7][25] = 4'h0;
    SS4[8][25] = 4'h0;
    SS4[9][25] = 4'h0;
    SS4[10][25] = 4'h0;
    SS4[11][25] = 4'h0;
    SS4[12][25] = 4'hE;
    SS4[13][25] = 4'hE;
    SS4[14][25] = 4'hE;
    SS4[15][25] = 4'hE;
    SS4[16][25] = 4'hE;
    SS4[17][25] = 4'hE;
    SS4[18][25] = 4'hD;
    SS4[19][25] = 4'hD;
    SS4[20][25] = 4'hD;
    SS4[21][25] = 4'hC;
    SS4[22][25] = 4'hC;
    SS4[23][25] = 4'hC;
    SS4[24][25] = 4'hD;
    SS4[25][25] = 4'hD;
    SS4[26][25] = 4'hD;
    SS4[27][25] = 4'hA;
    SS4[28][25] = 4'hA;
    SS4[29][25] = 4'hA;
    SS4[30][25] = 4'hC;
    SS4[31][25] = 4'hC;
    SS4[32][25] = 4'hC;
    SS4[33][25] = 4'hC;
    SS4[34][25] = 4'hC;
    SS4[35][25] = 4'hC;
    SS4[36][25] = 4'hC;
    SS4[37][25] = 4'hC;
    SS4[38][25] = 4'hC;
    SS4[39][25] = 4'hC;
    SS4[40][25] = 4'hC;
    SS4[41][25] = 4'hC;
    SS4[42][25] = 4'hC;
    SS4[43][25] = 4'hC;
    SS4[44][25] = 4'hC;
    SS4[45][25] = 4'hC;
    SS4[46][25] = 4'hC;
    SS4[47][25] = 4'hC;
    SS4[0][26] = 4'h0;
    SS4[1][26] = 4'h0;
    SS4[2][26] = 4'h0;
    SS4[3][26] = 4'h0;
    SS4[4][26] = 4'h0;
    SS4[5][26] = 4'h0;
    SS4[6][26] = 4'h0;
    SS4[7][26] = 4'h0;
    SS4[8][26] = 4'h0;
    SS4[9][26] = 4'h0;
    SS4[10][26] = 4'h0;
    SS4[11][26] = 4'h0;
    SS4[12][26] = 4'hE;
    SS4[13][26] = 4'hE;
    SS4[14][26] = 4'hE;
    SS4[15][26] = 4'hE;
    SS4[16][26] = 4'hE;
    SS4[17][26] = 4'hE;
    SS4[18][26] = 4'hD;
    SS4[19][26] = 4'hD;
    SS4[20][26] = 4'hD;
    SS4[21][26] = 4'hC;
    SS4[22][26] = 4'hC;
    SS4[23][26] = 4'hC;
    SS4[24][26] = 4'hD;
    SS4[25][26] = 4'hD;
    SS4[26][26] = 4'hD;
    SS4[27][26] = 4'hA;
    SS4[28][26] = 4'hA;
    SS4[29][26] = 4'hA;
    SS4[30][26] = 4'hC;
    SS4[31][26] = 4'hC;
    SS4[32][26] = 4'hC;
    SS4[33][26] = 4'hC;
    SS4[34][26] = 4'hC;
    SS4[35][26] = 4'hC;
    SS4[36][26] = 4'hC;
    SS4[37][26] = 4'hC;
    SS4[38][26] = 4'hC;
    SS4[39][26] = 4'hC;
    SS4[40][26] = 4'hC;
    SS4[41][26] = 4'hC;
    SS4[42][26] = 4'hC;
    SS4[43][26] = 4'hC;
    SS4[44][26] = 4'hC;
    SS4[45][26] = 4'hC;
    SS4[46][26] = 4'hC;
    SS4[47][26] = 4'hC;
    SS4[0][27] = 4'h0;
    SS4[1][27] = 4'h0;
    SS4[2][27] = 4'h0;
    SS4[3][27] = 4'h0;
    SS4[4][27] = 4'h0;
    SS4[5][27] = 4'h0;
    SS4[6][27] = 4'h0;
    SS4[7][27] = 4'h0;
    SS4[8][27] = 4'h0;
    SS4[9][27] = 4'hE;
    SS4[10][27] = 4'hE;
    SS4[11][27] = 4'hE;
    SS4[12][27] = 4'hD;
    SS4[13][27] = 4'hD;
    SS4[14][27] = 4'hD;
    SS4[15][27] = 4'hC;
    SS4[16][27] = 4'hC;
    SS4[17][27] = 4'hC;
    SS4[18][27] = 4'hC;
    SS4[19][27] = 4'hC;
    SS4[20][27] = 4'hC;
    SS4[21][27] = 4'hC;
    SS4[22][27] = 4'hC;
    SS4[23][27] = 4'hC;
    SS4[24][27] = 4'hC;
    SS4[25][27] = 4'hC;
    SS4[26][27] = 4'hC;
    SS4[27][27] = 4'hD;
    SS4[28][27] = 4'hD;
    SS4[29][27] = 4'hD;
    SS4[30][27] = 4'hC;
    SS4[31][27] = 4'hC;
    SS4[32][27] = 4'hC;
    SS4[33][27] = 4'hD;
    SS4[34][27] = 4'hD;
    SS4[35][27] = 4'hD;
    SS4[36][27] = 4'hD;
    SS4[37][27] = 4'hD;
    SS4[38][27] = 4'hD;
    SS4[39][27] = 4'hD;
    SS4[40][27] = 4'hD;
    SS4[41][27] = 4'hD;
    SS4[42][27] = 4'h0;
    SS4[43][27] = 4'h0;
    SS4[44][27] = 4'h0;
    SS4[45][27] = 4'h0;
    SS4[46][27] = 4'h0;
    SS4[47][27] = 4'h0;
    SS4[0][28] = 4'h0;
    SS4[1][28] = 4'h0;
    SS4[2][28] = 4'h0;
    SS4[3][28] = 4'h0;
    SS4[4][28] = 4'h0;
    SS4[5][28] = 4'h0;
    SS4[6][28] = 4'h0;
    SS4[7][28] = 4'h0;
    SS4[8][28] = 4'h0;
    SS4[9][28] = 4'hE;
    SS4[10][28] = 4'hE;
    SS4[11][28] = 4'hE;
    SS4[12][28] = 4'hD;
    SS4[13][28] = 4'hD;
    SS4[14][28] = 4'hD;
    SS4[15][28] = 4'hC;
    SS4[16][28] = 4'hC;
    SS4[17][28] = 4'hC;
    SS4[18][28] = 4'hC;
    SS4[19][28] = 4'hC;
    SS4[20][28] = 4'hC;
    SS4[21][28] = 4'hC;
    SS4[22][28] = 4'hC;
    SS4[23][28] = 4'hC;
    SS4[24][28] = 4'hC;
    SS4[25][28] = 4'hC;
    SS4[26][28] = 4'hC;
    SS4[27][28] = 4'hD;
    SS4[28][28] = 4'hD;
    SS4[29][28] = 4'hD;
    SS4[30][28] = 4'hC;
    SS4[31][28] = 4'hC;
    SS4[32][28] = 4'hC;
    SS4[33][28] = 4'hD;
    SS4[34][28] = 4'hD;
    SS4[35][28] = 4'hD;
    SS4[36][28] = 4'hD;
    SS4[37][28] = 4'hD;
    SS4[38][28] = 4'hD;
    SS4[39][28] = 4'hD;
    SS4[40][28] = 4'hD;
    SS4[41][28] = 4'hD;
    SS4[42][28] = 4'h0;
    SS4[43][28] = 4'h0;
    SS4[44][28] = 4'h0;
    SS4[45][28] = 4'h0;
    SS4[46][28] = 4'h0;
    SS4[47][28] = 4'h0;
    SS4[0][29] = 4'h0;
    SS4[1][29] = 4'h0;
    SS4[2][29] = 4'h0;
    SS4[3][29] = 4'h0;
    SS4[4][29] = 4'h0;
    SS4[5][29] = 4'h0;
    SS4[6][29] = 4'h0;
    SS4[7][29] = 4'h0;
    SS4[8][29] = 4'h0;
    SS4[9][29] = 4'hE;
    SS4[10][29] = 4'hE;
    SS4[11][29] = 4'hE;
    SS4[12][29] = 4'hD;
    SS4[13][29] = 4'hD;
    SS4[14][29] = 4'hD;
    SS4[15][29] = 4'hC;
    SS4[16][29] = 4'hC;
    SS4[17][29] = 4'hC;
    SS4[18][29] = 4'hC;
    SS4[19][29] = 4'hC;
    SS4[20][29] = 4'hC;
    SS4[21][29] = 4'hC;
    SS4[22][29] = 4'hC;
    SS4[23][29] = 4'hC;
    SS4[24][29] = 4'hC;
    SS4[25][29] = 4'hC;
    SS4[26][29] = 4'hC;
    SS4[27][29] = 4'hD;
    SS4[28][29] = 4'hD;
    SS4[29][29] = 4'hD;
    SS4[30][29] = 4'hC;
    SS4[31][29] = 4'hC;
    SS4[32][29] = 4'hC;
    SS4[33][29] = 4'hD;
    SS4[34][29] = 4'hD;
    SS4[35][29] = 4'hD;
    SS4[36][29] = 4'hD;
    SS4[37][29] = 4'hD;
    SS4[38][29] = 4'hD;
    SS4[39][29] = 4'hD;
    SS4[40][29] = 4'hD;
    SS4[41][29] = 4'hD;
    SS4[42][29] = 4'h0;
    SS4[43][29] = 4'h0;
    SS4[44][29] = 4'h0;
    SS4[45][29] = 4'h0;
    SS4[46][29] = 4'h0;
    SS4[47][29] = 4'h0;
    SS4[0][30] = 4'h0;
    SS4[1][30] = 4'h0;
    SS4[2][30] = 4'h0;
    SS4[3][30] = 4'h0;
    SS4[4][30] = 4'h0;
    SS4[5][30] = 4'h0;
    SS4[6][30] = 4'hE;
    SS4[7][30] = 4'hE;
    SS4[8][30] = 4'hE;
    SS4[9][30] = 4'hD;
    SS4[10][30] = 4'hD;
    SS4[11][30] = 4'hD;
    SS4[12][30] = 4'hC;
    SS4[13][30] = 4'hC;
    SS4[14][30] = 4'hC;
    SS4[15][30] = 4'hC;
    SS4[16][30] = 4'hC;
    SS4[17][30] = 4'hC;
    SS4[18][30] = 4'hC;
    SS4[19][30] = 4'hC;
    SS4[20][30] = 4'hC;
    SS4[21][30] = 4'hE;
    SS4[22][30] = 4'hE;
    SS4[23][30] = 4'hE;
    SS4[24][30] = 4'hD;
    SS4[25][30] = 4'hD;
    SS4[26][30] = 4'hD;
    SS4[27][30] = 4'hD;
    SS4[28][30] = 4'hD;
    SS4[29][30] = 4'hD;
    SS4[30][30] = 4'h0;
    SS4[31][30] = 4'h0;
    SS4[32][30] = 4'h0;
    SS4[33][30] = 4'h0;
    SS4[34][30] = 4'h0;
    SS4[35][30] = 4'h0;
    SS4[36][30] = 4'h0;
    SS4[37][30] = 4'h0;
    SS4[38][30] = 4'h0;
    SS4[39][30] = 4'h0;
    SS4[40][30] = 4'h0;
    SS4[41][30] = 4'h0;
    SS4[42][30] = 4'h0;
    SS4[43][30] = 4'h0;
    SS4[44][30] = 4'h0;
    SS4[45][30] = 4'h0;
    SS4[46][30] = 4'h0;
    SS4[47][30] = 4'h0;
    SS4[0][31] = 4'h0;
    SS4[1][31] = 4'h0;
    SS4[2][31] = 4'h0;
    SS4[3][31] = 4'h0;
    SS4[4][31] = 4'h0;
    SS4[5][31] = 4'h0;
    SS4[6][31] = 4'hE;
    SS4[7][31] = 4'hE;
    SS4[8][31] = 4'hE;
    SS4[9][31] = 4'hD;
    SS4[10][31] = 4'hD;
    SS4[11][31] = 4'hD;
    SS4[12][31] = 4'hC;
    SS4[13][31] = 4'hC;
    SS4[14][31] = 4'hC;
    SS4[15][31] = 4'hC;
    SS4[16][31] = 4'hC;
    SS4[17][31] = 4'hC;
    SS4[18][31] = 4'hC;
    SS4[19][31] = 4'hC;
    SS4[20][31] = 4'hC;
    SS4[21][31] = 4'hE;
    SS4[22][31] = 4'hE;
    SS4[23][31] = 4'hE;
    SS4[24][31] = 4'hD;
    SS4[25][31] = 4'hD;
    SS4[26][31] = 4'hD;
    SS4[27][31] = 4'hD;
    SS4[28][31] = 4'hD;
    SS4[29][31] = 4'hD;
    SS4[30][31] = 4'h0;
    SS4[31][31] = 4'h0;
    SS4[32][31] = 4'h0;
    SS4[33][31] = 4'h0;
    SS4[34][31] = 4'h0;
    SS4[35][31] = 4'h0;
    SS4[36][31] = 4'h0;
    SS4[37][31] = 4'h0;
    SS4[38][31] = 4'h0;
    SS4[39][31] = 4'h0;
    SS4[40][31] = 4'h0;
    SS4[41][31] = 4'h0;
    SS4[42][31] = 4'h0;
    SS4[43][31] = 4'h0;
    SS4[44][31] = 4'h0;
    SS4[45][31] = 4'h0;
    SS4[46][31] = 4'h0;
    SS4[47][31] = 4'h0;
    SS4[0][32] = 4'h0;
    SS4[1][32] = 4'h0;
    SS4[2][32] = 4'h0;
    SS4[3][32] = 4'h0;
    SS4[4][32] = 4'h0;
    SS4[5][32] = 4'h0;
    SS4[6][32] = 4'hE;
    SS4[7][32] = 4'hE;
    SS4[8][32] = 4'hE;
    SS4[9][32] = 4'hD;
    SS4[10][32] = 4'hD;
    SS4[11][32] = 4'hD;
    SS4[12][32] = 4'hC;
    SS4[13][32] = 4'hC;
    SS4[14][32] = 4'hC;
    SS4[15][32] = 4'hC;
    SS4[16][32] = 4'hC;
    SS4[17][32] = 4'hC;
    SS4[18][32] = 4'hC;
    SS4[19][32] = 4'hC;
    SS4[20][32] = 4'hC;
    SS4[21][32] = 4'hE;
    SS4[22][32] = 4'hE;
    SS4[23][32] = 4'hE;
    SS4[24][32] = 4'hD;
    SS4[25][32] = 4'hD;
    SS4[26][32] = 4'hD;
    SS4[27][32] = 4'hD;
    SS4[28][32] = 4'hD;
    SS4[29][32] = 4'hD;
    SS4[30][32] = 4'h0;
    SS4[31][32] = 4'h0;
    SS4[32][32] = 4'h0;
    SS4[33][32] = 4'h0;
    SS4[34][32] = 4'h0;
    SS4[35][32] = 4'h0;
    SS4[36][32] = 4'h0;
    SS4[37][32] = 4'h0;
    SS4[38][32] = 4'h0;
    SS4[39][32] = 4'h0;
    SS4[40][32] = 4'h0;
    SS4[41][32] = 4'h0;
    SS4[42][32] = 4'h0;
    SS4[43][32] = 4'h0;
    SS4[44][32] = 4'h0;
    SS4[45][32] = 4'h0;
    SS4[46][32] = 4'h0;
    SS4[47][32] = 4'h0;
    SS4[0][33] = 4'h0;
    SS4[1][33] = 4'h0;
    SS4[2][33] = 4'h0;
    SS4[3][33] = 4'hD;
    SS4[4][33] = 4'hD;
    SS4[5][33] = 4'hD;
    SS4[6][33] = 4'hC;
    SS4[7][33] = 4'hC;
    SS4[8][33] = 4'hC;
    SS4[9][33] = 4'hC;
    SS4[10][33] = 4'hC;
    SS4[11][33] = 4'hC;
    SS4[12][33] = 4'hC;
    SS4[13][33] = 4'hC;
    SS4[14][33] = 4'hC;
    SS4[15][33] = 4'hC;
    SS4[16][33] = 4'hC;
    SS4[17][33] = 4'hC;
    SS4[18][33] = 4'hE;
    SS4[19][33] = 4'hE;
    SS4[20][33] = 4'hE;
    SS4[21][33] = 4'hD;
    SS4[22][33] = 4'hD;
    SS4[23][33] = 4'hD;
    SS4[24][33] = 4'hD;
    SS4[25][33] = 4'hD;
    SS4[26][33] = 4'hD;
    SS4[27][33] = 4'h3;
    SS4[28][33] = 4'h3;
    SS4[29][33] = 4'h3;
    SS4[30][33] = 4'h0;
    SS4[31][33] = 4'h0;
    SS4[32][33] = 4'h0;
    SS4[33][33] = 4'h0;
    SS4[34][33] = 4'h0;
    SS4[35][33] = 4'h0;
    SS4[36][33] = 4'h0;
    SS4[37][33] = 4'h0;
    SS4[38][33] = 4'h0;
    SS4[39][33] = 4'h0;
    SS4[40][33] = 4'h0;
    SS4[41][33] = 4'h0;
    SS4[42][33] = 4'h0;
    SS4[43][33] = 4'h0;
    SS4[44][33] = 4'h0;
    SS4[45][33] = 4'h0;
    SS4[46][33] = 4'h0;
    SS4[47][33] = 4'h0;
    SS4[0][34] = 4'h0;
    SS4[1][34] = 4'h0;
    SS4[2][34] = 4'h0;
    SS4[3][34] = 4'hD;
    SS4[4][34] = 4'hD;
    SS4[5][34] = 4'hD;
    SS4[6][34] = 4'hC;
    SS4[7][34] = 4'hC;
    SS4[8][34] = 4'hC;
    SS4[9][34] = 4'hC;
    SS4[10][34] = 4'hC;
    SS4[11][34] = 4'hC;
    SS4[12][34] = 4'hC;
    SS4[13][34] = 4'hC;
    SS4[14][34] = 4'hC;
    SS4[15][34] = 4'hC;
    SS4[16][34] = 4'hC;
    SS4[17][34] = 4'hC;
    SS4[18][34] = 4'hE;
    SS4[19][34] = 4'hE;
    SS4[20][34] = 4'hE;
    SS4[21][34] = 4'hD;
    SS4[22][34] = 4'hD;
    SS4[23][34] = 4'hD;
    SS4[24][34] = 4'hD;
    SS4[25][34] = 4'hD;
    SS4[26][34] = 4'hD;
    SS4[27][34] = 4'h3;
    SS4[28][34] = 4'h3;
    SS4[29][34] = 4'h3;
    SS4[30][34] = 4'h0;
    SS4[31][34] = 4'h0;
    SS4[32][34] = 4'h0;
    SS4[33][34] = 4'h0;
    SS4[34][34] = 4'h0;
    SS4[35][34] = 4'h0;
    SS4[36][34] = 4'h0;
    SS4[37][34] = 4'h0;
    SS4[38][34] = 4'h0;
    SS4[39][34] = 4'h0;
    SS4[40][34] = 4'h0;
    SS4[41][34] = 4'h0;
    SS4[42][34] = 4'h0;
    SS4[43][34] = 4'h0;
    SS4[44][34] = 4'h0;
    SS4[45][34] = 4'h0;
    SS4[46][34] = 4'h0;
    SS4[47][34] = 4'h0;
    SS4[0][35] = 4'h0;
    SS4[1][35] = 4'h0;
    SS4[2][35] = 4'h0;
    SS4[3][35] = 4'hD;
    SS4[4][35] = 4'hD;
    SS4[5][35] = 4'hD;
    SS4[6][35] = 4'hC;
    SS4[7][35] = 4'hC;
    SS4[8][35] = 4'hC;
    SS4[9][35] = 4'hC;
    SS4[10][35] = 4'hC;
    SS4[11][35] = 4'hC;
    SS4[12][35] = 4'hC;
    SS4[13][35] = 4'hC;
    SS4[14][35] = 4'hC;
    SS4[15][35] = 4'hC;
    SS4[16][35] = 4'hC;
    SS4[17][35] = 4'hC;
    SS4[18][35] = 4'hE;
    SS4[19][35] = 4'hE;
    SS4[20][35] = 4'hE;
    SS4[21][35] = 4'hD;
    SS4[22][35] = 4'hD;
    SS4[23][35] = 4'hD;
    SS4[24][35] = 4'hD;
    SS4[25][35] = 4'hD;
    SS4[26][35] = 4'hD;
    SS4[27][35] = 4'h3;
    SS4[28][35] = 4'h3;
    SS4[29][35] = 4'h3;
    SS4[30][35] = 4'h0;
    SS4[31][35] = 4'h0;
    SS4[32][35] = 4'h0;
    SS4[33][35] = 4'h0;
    SS4[34][35] = 4'h0;
    SS4[35][35] = 4'h0;
    SS4[36][35] = 4'h0;
    SS4[37][35] = 4'h0;
    SS4[38][35] = 4'h0;
    SS4[39][35] = 4'h0;
    SS4[40][35] = 4'h0;
    SS4[41][35] = 4'h0;
    SS4[42][35] = 4'h0;
    SS4[43][35] = 4'h0;
    SS4[44][35] = 4'h0;
    SS4[45][35] = 4'h0;
    SS4[46][35] = 4'h0;
    SS4[47][35] = 4'h0;
    SS4[0][36] = 4'hD;
    SS4[1][36] = 4'hD;
    SS4[2][36] = 4'hD;
    SS4[3][36] = 4'hC;
    SS4[4][36] = 4'hC;
    SS4[5][36] = 4'hC;
    SS4[6][36] = 4'hC;
    SS4[7][36] = 4'hC;
    SS4[8][36] = 4'hC;
    SS4[9][36] = 4'h0;
    SS4[10][36] = 4'h0;
    SS4[11][36] = 4'h0;
    SS4[12][36] = 4'h0;
    SS4[13][36] = 4'h0;
    SS4[14][36] = 4'h0;
    SS4[15][36] = 4'hE;
    SS4[16][36] = 4'hE;
    SS4[17][36] = 4'hE;
    SS4[18][36] = 4'hE;
    SS4[19][36] = 4'hE;
    SS4[20][36] = 4'hE;
    SS4[21][36] = 4'hD;
    SS4[22][36] = 4'hD;
    SS4[23][36] = 4'hD;
    SS4[24][36] = 4'h0;
    SS4[25][36] = 4'h0;
    SS4[26][36] = 4'h0;
    SS4[27][36] = 4'h0;
    SS4[28][36] = 4'h0;
    SS4[29][36] = 4'h0;
    SS4[30][36] = 4'h0;
    SS4[31][36] = 4'h0;
    SS4[32][36] = 4'h0;
    SS4[33][36] = 4'h0;
    SS4[34][36] = 4'h0;
    SS4[35][36] = 4'h0;
    SS4[36][36] = 4'h0;
    SS4[37][36] = 4'h0;
    SS4[38][36] = 4'h0;
    SS4[39][36] = 4'h0;
    SS4[40][36] = 4'h0;
    SS4[41][36] = 4'h0;
    SS4[42][36] = 4'h0;
    SS4[43][36] = 4'h0;
    SS4[44][36] = 4'h0;
    SS4[45][36] = 4'h0;
    SS4[46][36] = 4'h0;
    SS4[47][36] = 4'h0;
    SS4[0][37] = 4'hD;
    SS4[1][37] = 4'hD;
    SS4[2][37] = 4'hD;
    SS4[3][37] = 4'hC;
    SS4[4][37] = 4'hC;
    SS4[5][37] = 4'hC;
    SS4[6][37] = 4'hC;
    SS4[7][37] = 4'hC;
    SS4[8][37] = 4'hC;
    SS4[9][37] = 4'h0;
    SS4[10][37] = 4'h0;
    SS4[11][37] = 4'h0;
    SS4[12][37] = 4'h0;
    SS4[13][37] = 4'h0;
    SS4[14][37] = 4'h0;
    SS4[15][37] = 4'hE;
    SS4[16][37] = 4'hE;
    SS4[17][37] = 4'hE;
    SS4[18][37] = 4'hE;
    SS4[19][37] = 4'hE;
    SS4[20][37] = 4'hE;
    SS4[21][37] = 4'hD;
    SS4[22][37] = 4'hD;
    SS4[23][37] = 4'hD;
    SS4[24][37] = 4'h0;
    SS4[25][37] = 4'h0;
    SS4[26][37] = 4'h0;
    SS4[27][37] = 4'h0;
    SS4[28][37] = 4'h0;
    SS4[29][37] = 4'h0;
    SS4[30][37] = 4'h0;
    SS4[31][37] = 4'h0;
    SS4[32][37] = 4'h0;
    SS4[33][37] = 4'h0;
    SS4[34][37] = 4'h0;
    SS4[35][37] = 4'h0;
    SS4[36][37] = 4'h0;
    SS4[37][37] = 4'h0;
    SS4[38][37] = 4'h0;
    SS4[39][37] = 4'h0;
    SS4[40][37] = 4'h0;
    SS4[41][37] = 4'h0;
    SS4[42][37] = 4'h0;
    SS4[43][37] = 4'h0;
    SS4[44][37] = 4'h0;
    SS4[45][37] = 4'h0;
    SS4[46][37] = 4'h0;
    SS4[47][37] = 4'h0;
    SS4[0][38] = 4'hD;
    SS4[1][38] = 4'hD;
    SS4[2][38] = 4'hD;
    SS4[3][38] = 4'hC;
    SS4[4][38] = 4'hC;
    SS4[5][38] = 4'hC;
    SS4[6][38] = 4'hC;
    SS4[7][38] = 4'hC;
    SS4[8][38] = 4'hC;
    SS4[9][38] = 4'h0;
    SS4[10][38] = 4'h0;
    SS4[11][38] = 4'h0;
    SS4[12][38] = 4'h0;
    SS4[13][38] = 4'h0;
    SS4[14][38] = 4'h0;
    SS4[15][38] = 4'hE;
    SS4[16][38] = 4'hE;
    SS4[17][38] = 4'hE;
    SS4[18][38] = 4'hE;
    SS4[19][38] = 4'hE;
    SS4[20][38] = 4'hE;
    SS4[21][38] = 4'hD;
    SS4[22][38] = 4'hD;
    SS4[23][38] = 4'hD;
    SS4[24][38] = 4'h0;
    SS4[25][38] = 4'h0;
    SS4[26][38] = 4'h0;
    SS4[27][38] = 4'h0;
    SS4[28][38] = 4'h0;
    SS4[29][38] = 4'h0;
    SS4[30][38] = 4'h0;
    SS4[31][38] = 4'h0;
    SS4[32][38] = 4'h0;
    SS4[33][38] = 4'h0;
    SS4[34][38] = 4'h0;
    SS4[35][38] = 4'h0;
    SS4[36][38] = 4'h0;
    SS4[37][38] = 4'h0;
    SS4[38][38] = 4'h0;
    SS4[39][38] = 4'h0;
    SS4[40][38] = 4'h0;
    SS4[41][38] = 4'h0;
    SS4[42][38] = 4'h0;
    SS4[43][38] = 4'h0;
    SS4[44][38] = 4'h0;
    SS4[45][38] = 4'h0;
    SS4[46][38] = 4'h0;
    SS4[47][38] = 4'h0;
    SS4[0][39] = 4'h0;
    SS4[1][39] = 4'h0;
    SS4[2][39] = 4'h0;
    SS4[3][39] = 4'h0;
    SS4[4][39] = 4'h0;
    SS4[5][39] = 4'h0;
    SS4[6][39] = 4'h0;
    SS4[7][39] = 4'h0;
    SS4[8][39] = 4'h0;
    SS4[9][39] = 4'h0;
    SS4[10][39] = 4'h0;
    SS4[11][39] = 4'h0;
    SS4[12][39] = 4'h0;
    SS4[13][39] = 4'h0;
    SS4[14][39] = 4'h0;
    SS4[15][39] = 4'hE;
    SS4[16][39] = 4'hE;
    SS4[17][39] = 4'hE;
    SS4[18][39] = 4'hD;
    SS4[19][39] = 4'hD;
    SS4[20][39] = 4'hD;
    SS4[21][39] = 4'h3;
    SS4[22][39] = 4'h3;
    SS4[23][39] = 4'h3;
    SS4[24][39] = 4'h0;
    SS4[25][39] = 4'h0;
    SS4[26][39] = 4'h0;
    SS4[27][39] = 4'h0;
    SS4[28][39] = 4'h0;
    SS4[29][39] = 4'h0;
    SS4[30][39] = 4'h0;
    SS4[31][39] = 4'h0;
    SS4[32][39] = 4'h0;
    SS4[33][39] = 4'h0;
    SS4[34][39] = 4'h0;
    SS4[35][39] = 4'h0;
    SS4[36][39] = 4'h0;
    SS4[37][39] = 4'h0;
    SS4[38][39] = 4'h0;
    SS4[39][39] = 4'h0;
    SS4[40][39] = 4'h0;
    SS4[41][39] = 4'h0;
    SS4[42][39] = 4'h0;
    SS4[43][39] = 4'h0;
    SS4[44][39] = 4'h0;
    SS4[45][39] = 4'h0;
    SS4[46][39] = 4'h0;
    SS4[47][39] = 4'h0;
    SS4[0][40] = 4'h0;
    SS4[1][40] = 4'h0;
    SS4[2][40] = 4'h0;
    SS4[3][40] = 4'h0;
    SS4[4][40] = 4'h0;
    SS4[5][40] = 4'h0;
    SS4[6][40] = 4'h0;
    SS4[7][40] = 4'h0;
    SS4[8][40] = 4'h0;
    SS4[9][40] = 4'h0;
    SS4[10][40] = 4'h0;
    SS4[11][40] = 4'h0;
    SS4[12][40] = 4'h0;
    SS4[13][40] = 4'h0;
    SS4[14][40] = 4'h0;
    SS4[15][40] = 4'hE;
    SS4[16][40] = 4'hE;
    SS4[17][40] = 4'hE;
    SS4[18][40] = 4'hD;
    SS4[19][40] = 4'hD;
    SS4[20][40] = 4'hD;
    SS4[21][40] = 4'h3;
    SS4[22][40] = 4'h3;
    SS4[23][40] = 4'h3;
    SS4[24][40] = 4'h0;
    SS4[25][40] = 4'h0;
    SS4[26][40] = 4'h0;
    SS4[27][40] = 4'h0;
    SS4[28][40] = 4'h0;
    SS4[29][40] = 4'h0;
    SS4[30][40] = 4'h0;
    SS4[31][40] = 4'h0;
    SS4[32][40] = 4'h0;
    SS4[33][40] = 4'h0;
    SS4[34][40] = 4'h0;
    SS4[35][40] = 4'h0;
    SS4[36][40] = 4'h0;
    SS4[37][40] = 4'h0;
    SS4[38][40] = 4'h0;
    SS4[39][40] = 4'h0;
    SS4[40][40] = 4'h0;
    SS4[41][40] = 4'h0;
    SS4[42][40] = 4'h0;
    SS4[43][40] = 4'h0;
    SS4[44][40] = 4'h0;
    SS4[45][40] = 4'h0;
    SS4[46][40] = 4'h0;
    SS4[47][40] = 4'h0;
    SS4[0][41] = 4'h0;
    SS4[1][41] = 4'h0;
    SS4[2][41] = 4'h0;
    SS4[3][41] = 4'h0;
    SS4[4][41] = 4'h0;
    SS4[5][41] = 4'h0;
    SS4[6][41] = 4'h0;
    SS4[7][41] = 4'h0;
    SS4[8][41] = 4'h0;
    SS4[9][41] = 4'h0;
    SS4[10][41] = 4'h0;
    SS4[11][41] = 4'h0;
    SS4[12][41] = 4'h0;
    SS4[13][41] = 4'h0;
    SS4[14][41] = 4'h0;
    SS4[15][41] = 4'hE;
    SS4[16][41] = 4'hE;
    SS4[17][41] = 4'hE;
    SS4[18][41] = 4'hD;
    SS4[19][41] = 4'hD;
    SS4[20][41] = 4'hD;
    SS4[21][41] = 4'h3;
    SS4[22][41] = 4'h3;
    SS4[23][41] = 4'h3;
    SS4[24][41] = 4'h0;
    SS4[25][41] = 4'h0;
    SS4[26][41] = 4'h0;
    SS4[27][41] = 4'h0;
    SS4[28][41] = 4'h0;
    SS4[29][41] = 4'h0;
    SS4[30][41] = 4'h0;
    SS4[31][41] = 4'h0;
    SS4[32][41] = 4'h0;
    SS4[33][41] = 4'h0;
    SS4[34][41] = 4'h0;
    SS4[35][41] = 4'h0;
    SS4[36][41] = 4'h0;
    SS4[37][41] = 4'h0;
    SS4[38][41] = 4'h0;
    SS4[39][41] = 4'h0;
    SS4[40][41] = 4'h0;
    SS4[41][41] = 4'h0;
    SS4[42][41] = 4'h0;
    SS4[43][41] = 4'h0;
    SS4[44][41] = 4'h0;
    SS4[45][41] = 4'h0;
    SS4[46][41] = 4'h0;
    SS4[47][41] = 4'h0;
    SS4[0][42] = 4'h0;
    SS4[1][42] = 4'h0;
    SS4[2][42] = 4'h0;
    SS4[3][42] = 4'h0;
    SS4[4][42] = 4'h0;
    SS4[5][42] = 4'h0;
    SS4[6][42] = 4'h0;
    SS4[7][42] = 4'h0;
    SS4[8][42] = 4'h0;
    SS4[9][42] = 4'h0;
    SS4[10][42] = 4'h0;
    SS4[11][42] = 4'h0;
    SS4[12][42] = 4'h0;
    SS4[13][42] = 4'h0;
    SS4[14][42] = 4'h0;
    SS4[15][42] = 4'hD;
    SS4[16][42] = 4'hD;
    SS4[17][42] = 4'hD;
    SS4[18][42] = 4'hD;
    SS4[19][42] = 4'hD;
    SS4[20][42] = 4'hD;
    SS4[21][42] = 4'h0;
    SS4[22][42] = 4'h0;
    SS4[23][42] = 4'h0;
    SS4[24][42] = 4'h0;
    SS4[25][42] = 4'h0;
    SS4[26][42] = 4'h0;
    SS4[27][42] = 4'h0;
    SS4[28][42] = 4'h0;
    SS4[29][42] = 4'h0;
    SS4[30][42] = 4'h0;
    SS4[31][42] = 4'h0;
    SS4[32][42] = 4'h0;
    SS4[33][42] = 4'h0;
    SS4[34][42] = 4'h0;
    SS4[35][42] = 4'h0;
    SS4[36][42] = 4'h0;
    SS4[37][42] = 4'h0;
    SS4[38][42] = 4'h0;
    SS4[39][42] = 4'h0;
    SS4[40][42] = 4'h0;
    SS4[41][42] = 4'h0;
    SS4[42][42] = 4'h0;
    SS4[43][42] = 4'h0;
    SS4[44][42] = 4'h0;
    SS4[45][42] = 4'h0;
    SS4[46][42] = 4'h0;
    SS4[47][42] = 4'h0;
    SS4[0][43] = 4'h0;
    SS4[1][43] = 4'h0;
    SS4[2][43] = 4'h0;
    SS4[3][43] = 4'h0;
    SS4[4][43] = 4'h0;
    SS4[5][43] = 4'h0;
    SS4[6][43] = 4'h0;
    SS4[7][43] = 4'h0;
    SS4[8][43] = 4'h0;
    SS4[9][43] = 4'h0;
    SS4[10][43] = 4'h0;
    SS4[11][43] = 4'h0;
    SS4[12][43] = 4'h0;
    SS4[13][43] = 4'h0;
    SS4[14][43] = 4'h0;
    SS4[15][43] = 4'hD;
    SS4[16][43] = 4'hD;
    SS4[17][43] = 4'hD;
    SS4[18][43] = 4'hD;
    SS4[19][43] = 4'hD;
    SS4[20][43] = 4'hD;
    SS4[21][43] = 4'h0;
    SS4[22][43] = 4'h0;
    SS4[23][43] = 4'h0;
    SS4[24][43] = 4'h0;
    SS4[25][43] = 4'h0;
    SS4[26][43] = 4'h0;
    SS4[27][43] = 4'h0;
    SS4[28][43] = 4'h0;
    SS4[29][43] = 4'h0;
    SS4[30][43] = 4'h0;
    SS4[31][43] = 4'h0;
    SS4[32][43] = 4'h0;
    SS4[33][43] = 4'h0;
    SS4[34][43] = 4'h0;
    SS4[35][43] = 4'h0;
    SS4[36][43] = 4'h0;
    SS4[37][43] = 4'h0;
    SS4[38][43] = 4'h0;
    SS4[39][43] = 4'h0;
    SS4[40][43] = 4'h0;
    SS4[41][43] = 4'h0;
    SS4[42][43] = 4'h0;
    SS4[43][43] = 4'h0;
    SS4[44][43] = 4'h0;
    SS4[45][43] = 4'h0;
    SS4[46][43] = 4'h0;
    SS4[47][43] = 4'h0;
    SS4[0][44] = 4'h0;
    SS4[1][44] = 4'h0;
    SS4[2][44] = 4'h0;
    SS4[3][44] = 4'h0;
    SS4[4][44] = 4'h0;
    SS4[5][44] = 4'h0;
    SS4[6][44] = 4'h0;
    SS4[7][44] = 4'h0;
    SS4[8][44] = 4'h0;
    SS4[9][44] = 4'h0;
    SS4[10][44] = 4'h0;
    SS4[11][44] = 4'h0;
    SS4[12][44] = 4'h0;
    SS4[13][44] = 4'h0;
    SS4[14][44] = 4'h0;
    SS4[15][44] = 4'hD;
    SS4[16][44] = 4'hD;
    SS4[17][44] = 4'hD;
    SS4[18][44] = 4'hD;
    SS4[19][44] = 4'hD;
    SS4[20][44] = 4'hD;
    SS4[21][44] = 4'h0;
    SS4[22][44] = 4'h0;
    SS4[23][44] = 4'h0;
    SS4[24][44] = 4'h0;
    SS4[25][44] = 4'h0;
    SS4[26][44] = 4'h0;
    SS4[27][44] = 4'h0;
    SS4[28][44] = 4'h0;
    SS4[29][44] = 4'h0;
    SS4[30][44] = 4'h0;
    SS4[31][44] = 4'h0;
    SS4[32][44] = 4'h0;
    SS4[33][44] = 4'h0;
    SS4[34][44] = 4'h0;
    SS4[35][44] = 4'h0;
    SS4[36][44] = 4'h0;
    SS4[37][44] = 4'h0;
    SS4[38][44] = 4'h0;
    SS4[39][44] = 4'h0;
    SS4[40][44] = 4'h0;
    SS4[41][44] = 4'h0;
    SS4[42][44] = 4'h0;
    SS4[43][44] = 4'h0;
    SS4[44][44] = 4'h0;
    SS4[45][44] = 4'h0;
    SS4[46][44] = 4'h0;
    SS4[47][44] = 4'h0;
    SS4[0][45] = 4'h0;
    SS4[1][45] = 4'h0;
    SS4[2][45] = 4'h0;
    SS4[3][45] = 4'h0;
    SS4[4][45] = 4'h0;
    SS4[5][45] = 4'h0;
    SS4[6][45] = 4'h0;
    SS4[7][45] = 4'h0;
    SS4[8][45] = 4'h0;
    SS4[9][45] = 4'h0;
    SS4[10][45] = 4'h0;
    SS4[11][45] = 4'h0;
    SS4[12][45] = 4'h0;
    SS4[13][45] = 4'h0;
    SS4[14][45] = 4'h0;
    SS4[15][45] = 4'hD;
    SS4[16][45] = 4'hD;
    SS4[17][45] = 4'hD;
    SS4[18][45] = 4'h0;
    SS4[19][45] = 4'h0;
    SS4[20][45] = 4'h0;
    SS4[21][45] = 4'h0;
    SS4[22][45] = 4'h0;
    SS4[23][45] = 4'h0;
    SS4[24][45] = 4'h0;
    SS4[25][45] = 4'h0;
    SS4[26][45] = 4'h0;
    SS4[27][45] = 4'h0;
    SS4[28][45] = 4'h0;
    SS4[29][45] = 4'h0;
    SS4[30][45] = 4'h0;
    SS4[31][45] = 4'h0;
    SS4[32][45] = 4'h0;
    SS4[33][45] = 4'h0;
    SS4[34][45] = 4'h0;
    SS4[35][45] = 4'h0;
    SS4[36][45] = 4'h0;
    SS4[37][45] = 4'h0;
    SS4[38][45] = 4'h0;
    SS4[39][45] = 4'h0;
    SS4[40][45] = 4'h0;
    SS4[41][45] = 4'h0;
    SS4[42][45] = 4'h0;
    SS4[43][45] = 4'h0;
    SS4[44][45] = 4'h0;
    SS4[45][45] = 4'h0;
    SS4[46][45] = 4'h0;
    SS4[47][45] = 4'h0;
    SS4[0][46] = 4'h0;
    SS4[1][46] = 4'h0;
    SS4[2][46] = 4'h0;
    SS4[3][46] = 4'h0;
    SS4[4][46] = 4'h0;
    SS4[5][46] = 4'h0;
    SS4[6][46] = 4'h0;
    SS4[7][46] = 4'h0;
    SS4[8][46] = 4'h0;
    SS4[9][46] = 4'h0;
    SS4[10][46] = 4'h0;
    SS4[11][46] = 4'h0;
    SS4[12][46] = 4'h0;
    SS4[13][46] = 4'h0;
    SS4[14][46] = 4'h0;
    SS4[15][46] = 4'hD;
    SS4[16][46] = 4'hD;
    SS4[17][46] = 4'hD;
    SS4[18][46] = 4'h0;
    SS4[19][46] = 4'h0;
    SS4[20][46] = 4'h0;
    SS4[21][46] = 4'h0;
    SS4[22][46] = 4'h0;
    SS4[23][46] = 4'h0;
    SS4[24][46] = 4'h0;
    SS4[25][46] = 4'h0;
    SS4[26][46] = 4'h0;
    SS4[27][46] = 4'h0;
    SS4[28][46] = 4'h0;
    SS4[29][46] = 4'h0;
    SS4[30][46] = 4'h0;
    SS4[31][46] = 4'h0;
    SS4[32][46] = 4'h0;
    SS4[33][46] = 4'h0;
    SS4[34][46] = 4'h0;
    SS4[35][46] = 4'h0;
    SS4[36][46] = 4'h0;
    SS4[37][46] = 4'h0;
    SS4[38][46] = 4'h0;
    SS4[39][46] = 4'h0;
    SS4[40][46] = 4'h0;
    SS4[41][46] = 4'h0;
    SS4[42][46] = 4'h0;
    SS4[43][46] = 4'h0;
    SS4[44][46] = 4'h0;
    SS4[45][46] = 4'h0;
    SS4[46][46] = 4'h0;
    SS4[47][46] = 4'h0;
    SS4[0][47] = 4'h0;
    SS4[1][47] = 4'h0;
    SS4[2][47] = 4'h0;
    SS4[3][47] = 4'h0;
    SS4[4][47] = 4'h0;
    SS4[5][47] = 4'h0;
    SS4[6][47] = 4'h0;
    SS4[7][47] = 4'h0;
    SS4[8][47] = 4'h0;
    SS4[9][47] = 4'h0;
    SS4[10][47] = 4'h0;
    SS4[11][47] = 4'h0;
    SS4[12][47] = 4'h0;
    SS4[13][47] = 4'h0;
    SS4[14][47] = 4'h0;
    SS4[15][47] = 4'hD;
    SS4[16][47] = 4'hD;
    SS4[17][47] = 4'hD;
    SS4[18][47] = 4'h0;
    SS4[19][47] = 4'h0;
    SS4[20][47] = 4'h0;
    SS4[21][47] = 4'h0;
    SS4[22][47] = 4'h0;
    SS4[23][47] = 4'h0;
    SS4[24][47] = 4'h0;
    SS4[25][47] = 4'h0;
    SS4[26][47] = 4'h0;
    SS4[27][47] = 4'h0;
    SS4[28][47] = 4'h0;
    SS4[29][47] = 4'h0;
    SS4[30][47] = 4'h0;
    SS4[31][47] = 4'h0;
    SS4[32][47] = 4'h0;
    SS4[33][47] = 4'h0;
    SS4[34][47] = 4'h0;
    SS4[35][47] = 4'h0;
    SS4[36][47] = 4'h0;
    SS4[37][47] = 4'h0;
    SS4[38][47] = 4'h0;
    SS4[39][47] = 4'h0;
    SS4[40][47] = 4'h0;
    SS4[41][47] = 4'h0;
    SS4[42][47] = 4'h0;
    SS4[43][47] = 4'h0;
    SS4[44][47] = 4'h0;
    SS4[45][47] = 4'h0;
    SS4[46][47] = 4'h0;
    SS4[47][47] = 4'h0;
 
//SS 5
    SS5[0][0] = 4'h0;
    SS5[1][0] = 4'h0;
    SS5[2][0] = 4'h0;
    SS5[3][0] = 4'h0;
    SS5[4][0] = 4'h0;
    SS5[5][0] = 4'h0;
    SS5[6][0] = 4'h0;
    SS5[7][0] = 4'h0;
    SS5[8][0] = 4'h0;
    SS5[9][0] = 4'h0;
    SS5[10][0] = 4'h0;
    SS5[11][0] = 4'h0;
    SS5[12][0] = 4'h0;
    SS5[13][0] = 4'h0;
    SS5[14][0] = 4'h0;
    SS5[15][0] = 4'h0;
    SS5[16][0] = 4'h0;
    SS5[17][0] = 4'h0;
    SS5[18][0] = 4'h0;
    SS5[19][0] = 4'h0;
    SS5[20][0] = 4'h0;
    SS5[21][0] = 4'h0;
    SS5[22][0] = 4'h0;
    SS5[23][0] = 4'h0;
    SS5[24][0] = 4'hD;
    SS5[25][0] = 4'hD;
    SS5[26][0] = 4'hD;
    SS5[27][0] = 4'h0;
    SS5[28][0] = 4'h0;
    SS5[29][0] = 4'h0;
    SS5[30][0] = 4'h0;
    SS5[31][0] = 4'h0;
    SS5[32][0] = 4'h0;
    SS5[33][0] = 4'h0;
    SS5[34][0] = 4'h0;
    SS5[35][0] = 4'h0;
    SS5[36][0] = 4'h0;
    SS5[37][0] = 4'h0;
    SS5[38][0] = 4'h0;
    SS5[39][0] = 4'h0;
    SS5[40][0] = 4'h0;
    SS5[41][0] = 4'h0;
    SS5[42][0] = 4'h0;
    SS5[43][0] = 4'h0;
    SS5[44][0] = 4'h0;
    SS5[45][0] = 4'h0;
    SS5[46][0] = 4'h0;
    SS5[47][0] = 4'h0;
    SS5[0][1] = 4'h0;
    SS5[1][1] = 4'h0;
    SS5[2][1] = 4'h0;
    SS5[3][1] = 4'h0;
    SS5[4][1] = 4'h0;
    SS5[5][1] = 4'h0;
    SS5[6][1] = 4'h0;
    SS5[7][1] = 4'h0;
    SS5[8][1] = 4'h0;
    SS5[9][1] = 4'h0;
    SS5[10][1] = 4'h0;
    SS5[11][1] = 4'h0;
    SS5[12][1] = 4'h0;
    SS5[13][1] = 4'h0;
    SS5[14][1] = 4'h0;
    SS5[15][1] = 4'h0;
    SS5[16][1] = 4'h0;
    SS5[17][1] = 4'h0;
    SS5[18][1] = 4'h0;
    SS5[19][1] = 4'h0;
    SS5[20][1] = 4'h0;
    SS5[21][1] = 4'h0;
    SS5[22][1] = 4'h0;
    SS5[23][1] = 4'h0;
    SS5[24][1] = 4'hD;
    SS5[25][1] = 4'hD;
    SS5[26][1] = 4'hD;
    SS5[27][1] = 4'h0;
    SS5[28][1] = 4'h0;
    SS5[29][1] = 4'h0;
    SS5[30][1] = 4'h0;
    SS5[31][1] = 4'h0;
    SS5[32][1] = 4'h0;
    SS5[33][1] = 4'h0;
    SS5[34][1] = 4'h0;
    SS5[35][1] = 4'h0;
    SS5[36][1] = 4'h0;
    SS5[37][1] = 4'h0;
    SS5[38][1] = 4'h0;
    SS5[39][1] = 4'h0;
    SS5[40][1] = 4'h0;
    SS5[41][1] = 4'h0;
    SS5[42][1] = 4'h0;
    SS5[43][1] = 4'h0;
    SS5[44][1] = 4'h0;
    SS5[45][1] = 4'h0;
    SS5[46][1] = 4'h0;
    SS5[47][1] = 4'h0;
    SS5[0][2] = 4'h0;
    SS5[1][2] = 4'h0;
    SS5[2][2] = 4'h0;
    SS5[3][2] = 4'h0;
    SS5[4][2] = 4'h0;
    SS5[5][2] = 4'h0;
    SS5[6][2] = 4'h0;
    SS5[7][2] = 4'hD;
    SS5[8][2] = 4'hD;
    SS5[9][2] = 4'hD;
    SS5[10][2] = 4'hC;
    SS5[11][2] = 4'h0;
    SS5[12][2] = 4'h0;
    SS5[13][2] = 4'h0;
    SS5[14][2] = 4'h0;
    SS5[15][2] = 4'h0;
    SS5[16][2] = 4'h0;
    SS5[17][2] = 4'h0;
    SS5[18][2] = 4'h0;
    SS5[19][2] = 4'h0;
    SS5[20][2] = 4'h0;
    SS5[21][2] = 4'h0;
    SS5[22][2] = 4'h0;
    SS5[23][2] = 4'hD;
    SS5[24][2] = 4'hD;
    SS5[25][2] = 4'hD;
    SS5[26][2] = 4'hE;
    SS5[27][2] = 4'h0;
    SS5[28][2] = 4'h0;
    SS5[29][2] = 4'h0;
    SS5[30][2] = 4'h0;
    SS5[31][2] = 4'h0;
    SS5[32][2] = 4'h0;
    SS5[33][2] = 4'h0;
    SS5[34][2] = 4'h0;
    SS5[35][2] = 4'h0;
    SS5[36][2] = 4'h0;
    SS5[37][2] = 4'h0;
    SS5[38][2] = 4'h0;
    SS5[39][2] = 4'h0;
    SS5[40][2] = 4'h0;
    SS5[41][2] = 4'h0;
    SS5[42][2] = 4'h0;
    SS5[43][2] = 4'h0;
    SS5[44][2] = 4'h0;
    SS5[45][2] = 4'h0;
    SS5[46][2] = 4'h0;
    SS5[47][2] = 4'h0;
    SS5[0][3] = 4'h0;
    SS5[1][3] = 4'h0;
    SS5[2][3] = 4'h0;
    SS5[3][3] = 4'h0;
    SS5[4][3] = 4'h0;
    SS5[5][3] = 4'h0;
    SS5[6][3] = 4'h0;
    SS5[7][3] = 4'hD;
    SS5[8][3] = 4'hD;
    SS5[9][3] = 4'hD;
    SS5[10][3] = 4'hC;
    SS5[11][3] = 4'hC;
    SS5[12][3] = 4'hC;
    SS5[13][3] = 4'h0;
    SS5[14][3] = 4'h0;
    SS5[15][3] = 4'h0;
    SS5[16][3] = 4'h0;
    SS5[17][3] = 4'h0;
    SS5[18][3] = 4'h0;
    SS5[19][3] = 4'h0;
    SS5[20][3] = 4'h0;
    SS5[21][3] = 4'h0;
    SS5[22][3] = 4'h0;
    SS5[23][3] = 4'hD;
    SS5[24][3] = 4'hD;
    SS5[25][3] = 4'hD;
    SS5[26][3] = 4'hD;
    SS5[27][3] = 4'hD;
    SS5[28][3] = 4'hD;
    SS5[29][3] = 4'h0;
    SS5[30][3] = 4'h0;
    SS5[31][3] = 4'h0;
    SS5[32][3] = 4'h0;
    SS5[33][3] = 4'h0;
    SS5[34][3] = 4'h0;
    SS5[35][3] = 4'h0;
    SS5[36][3] = 4'h0;
    SS5[37][3] = 4'h0;
    SS5[38][3] = 4'h0;
    SS5[39][3] = 4'h0;
    SS5[40][3] = 4'h0;
    SS5[41][3] = 4'h0;
    SS5[42][3] = 4'h0;
    SS5[43][3] = 4'h0;
    SS5[44][3] = 4'h0;
    SS5[45][3] = 4'h0;
    SS5[46][3] = 4'h0;
    SS5[47][3] = 4'h0;
    SS5[0][4] = 4'h0;
    SS5[1][4] = 4'h0;
    SS5[2][4] = 4'h0;
    SS5[3][4] = 4'h0;
    SS5[4][4] = 4'h0;
    SS5[5][4] = 4'h0;
    SS5[6][4] = 4'h0;
    SS5[7][4] = 4'h0;
    SS5[8][4] = 4'hD;
    SS5[9][4] = 4'hD;
    SS5[10][4] = 4'hC;
    SS5[11][4] = 4'hC;
    SS5[12][4] = 4'hC;
    SS5[13][4] = 4'hC;
    SS5[14][4] = 4'hC;
    SS5[15][4] = 4'hC;
    SS5[16][4] = 4'h0;
    SS5[17][4] = 4'h0;
    SS5[18][4] = 4'h0;
    SS5[19][4] = 4'h0;
    SS5[20][4] = 4'h0;
    SS5[21][4] = 4'h0;
    SS5[22][4] = 4'hE;
    SS5[23][4] = 4'hD;
    SS5[24][4] = 4'hD;
    SS5[25][4] = 4'hD;
    SS5[26][4] = 4'hD;
    SS5[27][4] = 4'hD;
    SS5[28][4] = 4'hD;
    SS5[29][4] = 4'h0;
    SS5[30][4] = 4'h0;
    SS5[31][4] = 4'h0;
    SS5[32][4] = 4'h0;
    SS5[33][4] = 4'h0;
    SS5[34][4] = 4'h0;
    SS5[35][4] = 4'h0;
    SS5[36][4] = 4'h0;
    SS5[37][4] = 4'h0;
    SS5[38][4] = 4'h0;
    SS5[39][4] = 4'h0;
    SS5[40][4] = 4'h0;
    SS5[41][4] = 4'h0;
    SS5[42][4] = 4'h0;
    SS5[43][4] = 4'h0;
    SS5[44][4] = 4'h0;
    SS5[45][4] = 4'h0;
    SS5[46][4] = 4'h0;
    SS5[47][4] = 4'h0;
    SS5[0][5] = 4'h0;
    SS5[1][5] = 4'h0;
    SS5[2][5] = 4'h0;
    SS5[3][5] = 4'h0;
    SS5[4][5] = 4'h0;
    SS5[5][5] = 4'h0;
    SS5[6][5] = 4'h0;
    SS5[7][5] = 4'h0;
    SS5[8][5] = 4'h0;
    SS5[9][5] = 4'hD;
    SS5[10][5] = 4'hC;
    SS5[11][5] = 4'hC;
    SS5[12][5] = 4'hC;
    SS5[13][5] = 4'hC;
    SS5[14][5] = 4'hC;
    SS5[15][5] = 4'hC;
    SS5[16][5] = 4'h0;
    SS5[17][5] = 4'h0;
    SS5[18][5] = 4'h0;
    SS5[19][5] = 4'h0;
    SS5[20][5] = 4'h0;
    SS5[21][5] = 4'h0;
    SS5[22][5] = 4'hE;
    SS5[23][5] = 4'hE;
    SS5[24][5] = 4'hE;
    SS5[25][5] = 4'hD;
    SS5[26][5] = 4'hD;
    SS5[27][5] = 4'hD;
    SS5[28][5] = 4'h0;
    SS5[29][5] = 4'h0;
    SS5[30][5] = 4'h0;
    SS5[31][5] = 4'h0;
    SS5[32][5] = 4'h0;
    SS5[33][5] = 4'h0;
    SS5[34][5] = 4'h0;
    SS5[35][5] = 4'h0;
    SS5[36][5] = 4'h0;
    SS5[37][5] = 4'h0;
    SS5[38][5] = 4'h0;
    SS5[39][5] = 4'h0;
    SS5[40][5] = 4'h0;
    SS5[41][5] = 4'h0;
    SS5[42][5] = 4'h0;
    SS5[43][5] = 4'h0;
    SS5[44][5] = 4'h0;
    SS5[45][5] = 4'h0;
    SS5[46][5] = 4'h0;
    SS5[47][5] = 4'h0;
    SS5[0][6] = 4'h0;
    SS5[1][6] = 4'h0;
    SS5[2][6] = 4'h0;
    SS5[3][6] = 4'h0;
    SS5[4][6] = 4'h0;
    SS5[5][6] = 4'h0;
    SS5[6][6] = 4'h0;
    SS5[7][6] = 4'h0;
    SS5[8][6] = 4'h0;
    SS5[9][6] = 4'hD;
    SS5[10][6] = 4'hD;
    SS5[11][6] = 4'hD;
    SS5[12][6] = 4'hC;
    SS5[13][6] = 4'hC;
    SS5[14][6] = 4'hC;
    SS5[15][6] = 4'h0;
    SS5[16][6] = 4'h0;
    SS5[17][6] = 4'h0;
    SS5[18][6] = 4'h0;
    SS5[19][6] = 4'h0;
    SS5[20][6] = 4'h0;
    SS5[21][6] = 4'h0;
    SS5[22][6] = 4'hE;
    SS5[23][6] = 4'hE;
    SS5[24][6] = 4'hE;
    SS5[25][6] = 4'hD;
    SS5[26][6] = 4'hD;
    SS5[27][6] = 4'hD;
    SS5[28][6] = 4'h0;
    SS5[29][6] = 4'h0;
    SS5[30][6] = 4'h0;
    SS5[31][6] = 4'h0;
    SS5[32][6] = 4'h0;
    SS5[33][6] = 4'h0;
    SS5[34][6] = 4'h0;
    SS5[35][6] = 4'h0;
    SS5[36][6] = 4'h0;
    SS5[37][6] = 4'h0;
    SS5[38][6] = 4'h0;
    SS5[39][6] = 4'h0;
    SS5[40][6] = 4'h0;
    SS5[41][6] = 4'h0;
    SS5[42][6] = 4'h0;
    SS5[43][6] = 4'h0;
    SS5[44][6] = 4'h0;
    SS5[45][6] = 4'h0;
    SS5[46][6] = 4'h0;
    SS5[47][6] = 4'h0;
    SS5[0][7] = 4'h0;
    SS5[1][7] = 4'h0;
    SS5[2][7] = 4'h0;
    SS5[3][7] = 4'h0;
    SS5[4][7] = 4'h0;
    SS5[5][7] = 4'h0;
    SS5[6][7] = 4'h0;
    SS5[7][7] = 4'h0;
    SS5[8][7] = 4'hD;
    SS5[9][7] = 4'hD;
    SS5[10][7] = 4'hD;
    SS5[11][7] = 4'hD;
    SS5[12][7] = 4'hC;
    SS5[13][7] = 4'hC;
    SS5[14][7] = 4'hC;
    SS5[15][7] = 4'h0;
    SS5[16][7] = 4'h0;
    SS5[17][7] = 4'h0;
    SS5[18][7] = 4'h0;
    SS5[19][7] = 4'h0;
    SS5[20][7] = 4'h0;
    SS5[21][7] = 4'hE;
    SS5[22][7] = 4'hE;
    SS5[23][7] = 4'hE;
    SS5[24][7] = 4'hD;
    SS5[25][7] = 4'hD;
    SS5[26][7] = 4'hD;
    SS5[27][7] = 4'hD;
    SS5[28][7] = 4'h3;
    SS5[29][7] = 4'h3;
    SS5[30][7] = 4'h3;
    SS5[31][7] = 4'h0;
    SS5[32][7] = 4'h0;
    SS5[33][7] = 4'h0;
    SS5[34][7] = 4'h0;
    SS5[35][7] = 4'h0;
    SS5[36][7] = 4'h0;
    SS5[37][7] = 4'h0;
    SS5[38][7] = 4'h0;
    SS5[39][7] = 4'h0;
    SS5[40][7] = 4'h0;
    SS5[41][7] = 4'h0;
    SS5[42][7] = 4'h0;
    SS5[43][7] = 4'h0;
    SS5[44][7] = 4'h0;
    SS5[45][7] = 4'h0;
    SS5[46][7] = 4'h0;
    SS5[47][7] = 4'h0;
    SS5[0][8] = 4'h0;
    SS5[1][8] = 4'h0;
    SS5[2][8] = 4'h0;
    SS5[3][8] = 4'h0;
    SS5[4][8] = 4'h0;
    SS5[5][8] = 4'h0;
    SS5[6][8] = 4'h0;
    SS5[7][8] = 4'h0;
    SS5[8][8] = 4'h0;
    SS5[9][8] = 4'h0;
    SS5[10][8] = 4'hD;
    SS5[11][8] = 4'hC;
    SS5[12][8] = 4'hC;
    SS5[13][8] = 4'hC;
    SS5[14][8] = 4'hC;
    SS5[15][8] = 4'hC;
    SS5[16][8] = 4'hC;
    SS5[17][8] = 4'hC;
    SS5[18][8] = 4'h0;
    SS5[19][8] = 4'h0;
    SS5[20][8] = 4'h0;
    SS5[21][8] = 4'hE;
    SS5[22][8] = 4'hE;
    SS5[23][8] = 4'hE;
    SS5[24][8] = 4'hE;
    SS5[25][8] = 4'hD;
    SS5[26][8] = 4'hD;
    SS5[27][8] = 4'h3;
    SS5[28][8] = 4'h3;
    SS5[29][8] = 4'h3;
    SS5[30][8] = 4'h0;
    SS5[31][8] = 4'h0;
    SS5[32][8] = 4'h0;
    SS5[33][8] = 4'h0;
    SS5[34][8] = 4'h0;
    SS5[35][8] = 4'h0;
    SS5[36][8] = 4'h0;
    SS5[37][8] = 4'h0;
    SS5[38][8] = 4'h0;
    SS5[39][8] = 4'h0;
    SS5[40][8] = 4'h0;
    SS5[41][8] = 4'h0;
    SS5[42][8] = 4'h0;
    SS5[43][8] = 4'h0;
    SS5[44][8] = 4'h0;
    SS5[45][8] = 4'h0;
    SS5[46][8] = 4'h0;
    SS5[47][8] = 4'h0;
    SS5[0][9] = 4'h0;
    SS5[1][9] = 4'h0;
    SS5[2][9] = 4'h0;
    SS5[3][9] = 4'h0;
    SS5[4][9] = 4'h0;
    SS5[5][9] = 4'h0;
    SS5[6][9] = 4'h0;
    SS5[7][9] = 4'h0;
    SS5[8][9] = 4'h0;
    SS5[9][9] = 4'h0;
    SS5[10][9] = 4'h0;
    SS5[11][9] = 4'hE;
    SS5[12][9] = 4'hC;
    SS5[13][9] = 4'hC;
    SS5[14][9] = 4'hC;
    SS5[15][9] = 4'hC;
    SS5[16][9] = 4'hC;
    SS5[17][9] = 4'hC;
    SS5[18][9] = 4'hC;
    SS5[19][9] = 4'hC;
    SS5[20][9] = 4'hE;
    SS5[21][9] = 4'hE;
    SS5[22][9] = 4'hE;
    SS5[23][9] = 4'hE;
    SS5[24][9] = 4'hE;
    SS5[25][9] = 4'hE;
    SS5[26][9] = 4'hE;
    SS5[27][9] = 4'hD;
    SS5[28][9] = 4'h3;
    SS5[29][9] = 4'h3;
    SS5[30][9] = 4'h0;
    SS5[31][9] = 4'h0;
    SS5[32][9] = 4'h0;
    SS5[33][9] = 4'h0;
    SS5[34][9] = 4'h0;
    SS5[35][9] = 4'h0;
    SS5[36][9] = 4'h0;
    SS5[37][9] = 4'h0;
    SS5[38][9] = 4'h0;
    SS5[39][9] = 4'h0;
    SS5[40][9] = 4'h0;
    SS5[41][9] = 4'h0;
    SS5[42][9] = 4'h0;
    SS5[43][9] = 4'h0;
    SS5[44][9] = 4'h0;
    SS5[45][9] = 4'h0;
    SS5[46][9] = 4'h0;
    SS5[47][9] = 4'h0;
    SS5[0][10] = 4'h0;
    SS5[1][10] = 4'h0;
    SS5[2][10] = 4'h0;
    SS5[3][10] = 4'h0;
    SS5[4][10] = 4'h0;
    SS5[5][10] = 4'h0;
    SS5[6][10] = 4'h0;
    SS5[7][10] = 4'h0;
    SS5[8][10] = 4'h0;
    SS5[9][10] = 4'h0;
    SS5[10][10] = 4'hE;
    SS5[11][10] = 4'hE;
    SS5[12][10] = 4'hE;
    SS5[13][10] = 4'hE;
    SS5[14][10] = 4'hD;
    SS5[15][10] = 4'hC;
    SS5[16][10] = 4'hC;
    SS5[17][10] = 4'hC;
    SS5[18][10] = 4'hC;
    SS5[19][10] = 4'hC;
    SS5[20][10] = 4'hC;
    SS5[21][10] = 4'hC;
    SS5[22][10] = 4'hE;
    SS5[23][10] = 4'hE;
    SS5[24][10] = 4'hE;
    SS5[25][10] = 4'hE;
    SS5[26][10] = 4'hD;
    SS5[27][10] = 4'hD;
    SS5[28][10] = 4'hD;
    SS5[29][10] = 4'hD;
    SS5[30][10] = 4'h0;
    SS5[31][10] = 4'h0;
    SS5[32][10] = 4'h0;
    SS5[33][10] = 4'h0;
    SS5[34][10] = 4'h0;
    SS5[35][10] = 4'h0;
    SS5[36][10] = 4'h0;
    SS5[37][10] = 4'h0;
    SS5[38][10] = 4'h0;
    SS5[39][10] = 4'h0;
    SS5[40][10] = 4'h0;
    SS5[41][10] = 4'h0;
    SS5[42][10] = 4'h0;
    SS5[43][10] = 4'h0;
    SS5[44][10] = 4'h0;
    SS5[45][10] = 4'h0;
    SS5[46][10] = 4'h0;
    SS5[47][10] = 4'h0;
    SS5[0][11] = 4'h0;
    SS5[1][11] = 4'h0;
    SS5[2][11] = 4'h0;
    SS5[3][11] = 4'h0;
    SS5[4][11] = 4'h0;
    SS5[5][11] = 4'h0;
    SS5[6][11] = 4'h0;
    SS5[7][11] = 4'h0;
    SS5[8][11] = 4'h0;
    SS5[9][11] = 4'h0;
    SS5[10][11] = 4'hE;
    SS5[11][11] = 4'hE;
    SS5[12][11] = 4'hE;
    SS5[13][11] = 4'hD;
    SS5[14][11] = 4'hD;
    SS5[15][11] = 4'hD;
    SS5[16][11] = 4'hC;
    SS5[17][11] = 4'hC;
    SS5[18][11] = 4'hC;
    SS5[19][11] = 4'hC;
    SS5[20][11] = 4'hC;
    SS5[21][11] = 4'hC;
    SS5[22][11] = 4'hC;
    SS5[23][11] = 4'hE;
    SS5[24][11] = 4'hE;
    SS5[25][11] = 4'hE;
    SS5[26][11] = 4'hD;
    SS5[27][11] = 4'hD;
    SS5[28][11] = 4'hD;
    SS5[29][11] = 4'h0;
    SS5[30][11] = 4'h0;
    SS5[31][11] = 4'h0;
    SS5[32][11] = 4'h0;
    SS5[33][11] = 4'h0;
    SS5[34][11] = 4'h0;
    SS5[35][11] = 4'h0;
    SS5[36][11] = 4'h0;
    SS5[37][11] = 4'h0;
    SS5[38][11] = 4'h0;
    SS5[39][11] = 4'h0;
    SS5[40][11] = 4'h0;
    SS5[41][11] = 4'h0;
    SS5[42][11] = 4'h0;
    SS5[43][11] = 4'h0;
    SS5[44][11] = 4'h0;
    SS5[45][11] = 4'h0;
    SS5[46][11] = 4'h0;
    SS5[47][11] = 4'h0;
    SS5[0][12] = 4'h0;
    SS5[1][12] = 4'h0;
    SS5[2][12] = 4'h0;
    SS5[3][12] = 4'h0;
    SS5[4][12] = 4'h0;
    SS5[5][12] = 4'h0;
    SS5[6][12] = 4'h0;
    SS5[7][12] = 4'h0;
    SS5[8][12] = 4'h0;
    SS5[9][12] = 4'h0;
    SS5[10][12] = 4'h0;
    SS5[11][12] = 4'h0;
    SS5[12][12] = 4'hE;
    SS5[13][12] = 4'hD;
    SS5[14][12] = 4'hD;
    SS5[15][12] = 4'hD;
    SS5[16][12] = 4'hC;
    SS5[17][12] = 4'hC;
    SS5[18][12] = 4'hC;
    SS5[19][12] = 4'hC;
    SS5[20][12] = 4'hC;
    SS5[21][12] = 4'hC;
    SS5[22][12] = 4'hE;
    SS5[23][12] = 4'hE;
    SS5[24][12] = 4'hE;
    SS5[25][12] = 4'hE;
    SS5[26][12] = 4'hD;
    SS5[27][12] = 4'hD;
    SS5[28][12] = 4'hD;
    SS5[29][12] = 4'h0;
    SS5[30][12] = 4'h0;
    SS5[31][12] = 4'h0;
    SS5[32][12] = 4'h0;
    SS5[33][12] = 4'h0;
    SS5[34][12] = 4'h0;
    SS5[35][12] = 4'h0;
    SS5[36][12] = 4'h0;
    SS5[37][12] = 4'h0;
    SS5[38][12] = 4'h0;
    SS5[39][12] = 4'h0;
    SS5[40][12] = 4'h0;
    SS5[41][12] = 4'h0;
    SS5[42][12] = 4'h0;
    SS5[43][12] = 4'h0;
    SS5[44][12] = 4'h0;
    SS5[45][12] = 4'h0;
    SS5[46][12] = 4'h0;
    SS5[47][12] = 4'h0;
    SS5[0][13] = 4'h0;
    SS5[1][13] = 4'h0;
    SS5[2][13] = 4'h0;
    SS5[3][13] = 4'h0;
    SS5[4][13] = 4'h0;
    SS5[5][13] = 4'h0;
    SS5[6][13] = 4'h0;
    SS5[7][13] = 4'h0;
    SS5[8][13] = 4'h0;
    SS5[9][13] = 4'h0;
    SS5[10][13] = 4'h0;
    SS5[11][13] = 4'h0;
    SS5[12][13] = 4'hE;
    SS5[13][13] = 4'hE;
    SS5[14][13] = 4'hD;
    SS5[15][13] = 4'hD;
    SS5[16][13] = 4'hC;
    SS5[17][13] = 4'hC;
    SS5[18][13] = 4'hC;
    SS5[19][13] = 4'hC;
    SS5[20][13] = 4'hC;
    SS5[21][13] = 4'hC;
    SS5[22][13] = 4'hE;
    SS5[23][13] = 4'hE;
    SS5[24][13] = 4'hE;
    SS5[25][13] = 4'hD;
    SS5[26][13] = 4'hD;
    SS5[27][13] = 4'hD;
    SS5[28][13] = 4'hD;
    SS5[29][13] = 4'hD;
    SS5[30][13] = 4'h0;
    SS5[31][13] = 4'h0;
    SS5[32][13] = 4'h0;
    SS5[33][13] = 4'h0;
    SS5[34][13] = 4'h0;
    SS5[35][13] = 4'h0;
    SS5[36][13] = 4'h0;
    SS5[37][13] = 4'h0;
    SS5[38][13] = 4'h0;
    SS5[39][13] = 4'h0;
    SS5[40][13] = 4'h0;
    SS5[41][13] = 4'h0;
    SS5[42][13] = 4'h0;
    SS5[43][13] = 4'h0;
    SS5[44][13] = 4'h0;
    SS5[45][13] = 4'h0;
    SS5[46][13] = 4'h0;
    SS5[47][13] = 4'h0;
    SS5[0][14] = 4'h0;
    SS5[1][14] = 4'h0;
    SS5[2][14] = 4'h0;
    SS5[3][14] = 4'h0;
    SS5[4][14] = 4'h0;
    SS5[5][14] = 4'h0;
    SS5[6][14] = 4'h0;
    SS5[7][14] = 4'h0;
    SS5[8][14] = 4'h0;
    SS5[9][14] = 4'h0;
    SS5[10][14] = 4'h0;
    SS5[11][14] = 4'h0;
    SS5[12][14] = 4'hE;
    SS5[13][14] = 4'hE;
    SS5[14][14] = 4'hE;
    SS5[15][14] = 4'hD;
    SS5[16][14] = 4'hD;
    SS5[17][14] = 4'hC;
    SS5[18][14] = 4'hC;
    SS5[19][14] = 4'hC;
    SS5[20][14] = 4'hC;
    SS5[21][14] = 4'hC;
    SS5[22][14] = 4'hC;
    SS5[23][14] = 4'hC;
    SS5[24][14] = 4'hE;
    SS5[25][14] = 4'hD;
    SS5[26][14] = 4'hD;
    SS5[27][14] = 4'hD;
    SS5[28][14] = 4'hD;
    SS5[29][14] = 4'hD;
    SS5[30][14] = 4'hD;
    SS5[31][14] = 4'h3;
    SS5[32][14] = 4'h0;
    SS5[33][14] = 4'h0;
    SS5[34][14] = 4'h0;
    SS5[35][14] = 4'h0;
    SS5[36][14] = 4'h0;
    SS5[37][14] = 4'h0;
    SS5[38][14] = 4'h0;
    SS5[39][14] = 4'h0;
    SS5[40][14] = 4'h0;
    SS5[41][14] = 4'h0;
    SS5[42][14] = 4'h0;
    SS5[43][14] = 4'h0;
    SS5[44][14] = 4'h0;
    SS5[45][14] = 4'h0;
    SS5[46][14] = 4'h0;
    SS5[47][14] = 4'h0;
    SS5[0][15] = 4'h0;
    SS5[1][15] = 4'h0;
    SS5[2][15] = 4'h0;
    SS5[3][15] = 4'h0;
    SS5[4][15] = 4'h0;
    SS5[5][15] = 4'h0;
    SS5[6][15] = 4'h0;
    SS5[7][15] = 4'h0;
    SS5[8][15] = 4'h0;
    SS5[9][15] = 4'h0;
    SS5[10][15] = 4'h0;
    SS5[11][15] = 4'hE;
    SS5[12][15] = 4'hE;
    SS5[13][15] = 4'hE;
    SS5[14][15] = 4'hE;
    SS5[15][15] = 4'hD;
    SS5[16][15] = 4'hD;
    SS5[17][15] = 4'hD;
    SS5[18][15] = 4'hC;
    SS5[19][15] = 4'hC;
    SS5[20][15] = 4'hC;
    SS5[21][15] = 4'hC;
    SS5[22][15] = 4'hC;
    SS5[23][15] = 4'hC;
    SS5[24][15] = 4'hE;
    SS5[25][15] = 4'hE;
    SS5[26][15] = 4'hE;
    SS5[27][15] = 4'hD;
    SS5[28][15] = 4'hD;
    SS5[29][15] = 4'hD;
    SS5[30][15] = 4'hD;
    SS5[31][15] = 4'h3;
    SS5[32][15] = 4'h3;
    SS5[33][15] = 4'h3;
    SS5[34][15] = 4'h0;
    SS5[35][15] = 4'h0;
    SS5[36][15] = 4'h0;
    SS5[37][15] = 4'h0;
    SS5[38][15] = 4'h0;
    SS5[39][15] = 4'h0;
    SS5[40][15] = 4'h0;
    SS5[41][15] = 4'h0;
    SS5[42][15] = 4'h0;
    SS5[43][15] = 4'h0;
    SS5[44][15] = 4'h0;
    SS5[45][15] = 4'h0;
    SS5[46][15] = 4'h0;
    SS5[47][15] = 4'h0;
    SS5[0][16] = 4'h0;
    SS5[1][16] = 4'h0;
    SS5[2][16] = 4'h0;
    SS5[3][16] = 4'h0;
    SS5[4][16] = 4'h0;
    SS5[5][16] = 4'h0;
    SS5[6][16] = 4'h0;
    SS5[7][16] = 4'h0;
    SS5[8][16] = 4'h0;
    SS5[9][16] = 4'h0;
    SS5[10][16] = 4'h0;
    SS5[11][16] = 4'h0;
    SS5[12][16] = 4'h0;
    SS5[13][16] = 4'h0;
    SS5[14][16] = 4'hD;
    SS5[15][16] = 4'hD;
    SS5[16][16] = 4'hD;
    SS5[17][16] = 4'hC;
    SS5[18][16] = 4'hC;
    SS5[19][16] = 4'hC;
    SS5[20][16] = 4'hC;
    SS5[21][16] = 4'hC;
    SS5[22][16] = 4'hC;
    SS5[23][16] = 4'hC;
    SS5[24][16] = 4'hE;
    SS5[25][16] = 4'hE;
    SS5[26][16] = 4'hE;
    SS5[27][16] = 4'hD;
    SS5[28][16] = 4'hD;
    SS5[29][16] = 4'hD;
    SS5[30][16] = 4'h3;
    SS5[31][16] = 4'h3;
    SS5[32][16] = 4'h3;
    SS5[33][16] = 4'h3;
    SS5[34][16] = 4'h0;
    SS5[35][16] = 4'h0;
    SS5[36][16] = 4'h0;
    SS5[37][16] = 4'h0;
    SS5[38][16] = 4'h0;
    SS5[39][16] = 4'h0;
    SS5[40][16] = 4'h0;
    SS5[41][16] = 4'h0;
    SS5[42][16] = 4'h0;
    SS5[43][16] = 4'h0;
    SS5[44][16] = 4'h0;
    SS5[45][16] = 4'h0;
    SS5[46][16] = 4'h0;
    SS5[47][16] = 4'h0;
    SS5[0][17] = 4'h0;
    SS5[1][17] = 4'h0;
    SS5[2][17] = 4'h0;
    SS5[3][17] = 4'h0;
    SS5[4][17] = 4'h0;
    SS5[5][17] = 4'h0;
    SS5[6][17] = 4'h0;
    SS5[7][17] = 4'h0;
    SS5[8][17] = 4'h0;
    SS5[9][17] = 4'h0;
    SS5[10][17] = 4'h0;
    SS5[11][17] = 4'h0;
    SS5[12][17] = 4'h0;
    SS5[13][17] = 4'h0;
    SS5[14][17] = 4'hE;
    SS5[15][17] = 4'hE;
    SS5[16][17] = 4'hD;
    SS5[17][17] = 4'hC;
    SS5[18][17] = 4'hC;
    SS5[19][17] = 4'hC;
    SS5[20][17] = 4'hC;
    SS5[21][17] = 4'hC;
    SS5[22][17] = 4'hC;
    SS5[23][17] = 4'hC;
    SS5[24][17] = 4'hE;
    SS5[25][17] = 4'hE;
    SS5[26][17] = 4'hE;
    SS5[27][17] = 4'hD;
    SS5[28][17] = 4'hD;
    SS5[29][17] = 4'hD;
    SS5[30][17] = 4'hD;
    SS5[31][17] = 4'hD;
    SS5[32][17] = 4'h3;
    SS5[33][17] = 4'h0;
    SS5[34][17] = 4'h0;
    SS5[35][17] = 4'h0;
    SS5[36][17] = 4'h0;
    SS5[37][17] = 4'h0;
    SS5[38][17] = 4'h0;
    SS5[39][17] = 4'h0;
    SS5[40][17] = 4'h0;
    SS5[41][17] = 4'h0;
    SS5[42][17] = 4'h0;
    SS5[43][17] = 4'h0;
    SS5[44][17] = 4'h0;
    SS5[45][17] = 4'h0;
    SS5[46][17] = 4'h0;
    SS5[47][17] = 4'h0;
    SS5[0][18] = 4'h0;
    SS5[1][18] = 4'h0;
    SS5[2][18] = 4'h0;
    SS5[3][18] = 4'h0;
    SS5[4][18] = 4'h0;
    SS5[5][18] = 4'h0;
    SS5[6][18] = 4'h0;
    SS5[7][18] = 4'h0;
    SS5[8][18] = 4'h0;
    SS5[9][18] = 4'h0;
    SS5[10][18] = 4'h0;
    SS5[11][18] = 4'h0;
    SS5[12][18] = 4'h0;
    SS5[13][18] = 4'hE;
    SS5[14][18] = 4'hE;
    SS5[15][18] = 4'hE;
    SS5[16][18] = 4'hE;
    SS5[17][18] = 4'hE;
    SS5[18][18] = 4'hC;
    SS5[19][18] = 4'hC;
    SS5[20][18] = 4'hC;
    SS5[21][18] = 4'hC;
    SS5[22][18] = 4'hC;
    SS5[23][18] = 4'hC;
    SS5[24][18] = 4'hC;
    SS5[25][18] = 4'hC;
    SS5[26][18] = 4'hD;
    SS5[27][18] = 4'hD;
    SS5[28][18] = 4'hD;
    SS5[29][18] = 4'hD;
    SS5[30][18] = 4'hD;
    SS5[31][18] = 4'hD;
    SS5[32][18] = 4'hD;
    SS5[33][18] = 4'h0;
    SS5[34][18] = 4'h0;
    SS5[35][18] = 4'h0;
    SS5[36][18] = 4'h0;
    SS5[37][18] = 4'h0;
    SS5[38][18] = 4'h0;
    SS5[39][18] = 4'h0;
    SS5[40][18] = 4'h0;
    SS5[41][18] = 4'h0;
    SS5[42][18] = 4'h0;
    SS5[43][18] = 4'h0;
    SS5[44][18] = 4'h0;
    SS5[45][18] = 4'h0;
    SS5[46][18] = 4'h0;
    SS5[47][18] = 4'h0;
    SS5[0][19] = 4'h0;
    SS5[1][19] = 4'h0;
    SS5[2][19] = 4'h0;
    SS5[3][19] = 4'h0;
    SS5[4][19] = 4'h0;
    SS5[5][19] = 4'h0;
    SS5[6][19] = 4'h0;
    SS5[7][19] = 4'h0;
    SS5[8][19] = 4'h0;
    SS5[9][19] = 4'h0;
    SS5[10][19] = 4'h0;
    SS5[11][19] = 4'h0;
    SS5[12][19] = 4'h0;
    SS5[13][19] = 4'hE;
    SS5[14][19] = 4'hE;
    SS5[15][19] = 4'hE;
    SS5[16][19] = 4'hE;
    SS5[17][19] = 4'hE;
    SS5[18][19] = 4'hE;
    SS5[19][19] = 4'hD;
    SS5[20][19] = 4'hD;
    SS5[21][19] = 4'hC;
    SS5[22][19] = 4'hC;
    SS5[23][19] = 4'hC;
    SS5[24][19] = 4'hC;
    SS5[25][19] = 4'hC;
    SS5[26][19] = 4'hC;
    SS5[27][19] = 4'hC;
    SS5[28][19] = 4'hC;
    SS5[29][19] = 4'hD;
    SS5[30][19] = 4'hD;
    SS5[31][19] = 4'hD;
    SS5[32][19] = 4'h0;
    SS5[33][19] = 4'h0;
    SS5[34][19] = 4'h0;
    SS5[35][19] = 4'h0;
    SS5[36][19] = 4'h0;
    SS5[37][19] = 4'h0;
    SS5[38][19] = 4'h0;
    SS5[39][19] = 4'h0;
    SS5[40][19] = 4'h0;
    SS5[41][19] = 4'h0;
    SS5[42][19] = 4'h0;
    SS5[43][19] = 4'h0;
    SS5[44][19] = 4'h0;
    SS5[45][19] = 4'h0;
    SS5[46][19] = 4'h0;
    SS5[47][19] = 4'h0;
    SS5[0][20] = 4'h0;
    SS5[1][20] = 4'h0;
    SS5[2][20] = 4'h0;
    SS5[3][20] = 4'h0;
    SS5[4][20] = 4'h0;
    SS5[5][20] = 4'h0;
    SS5[6][20] = 4'h0;
    SS5[7][20] = 4'h0;
    SS5[8][20] = 4'h0;
    SS5[9][20] = 4'h0;
    SS5[10][20] = 4'h0;
    SS5[11][20] = 4'h0;
    SS5[12][20] = 4'h0;
    SS5[13][20] = 4'hE;
    SS5[14][20] = 4'hE;
    SS5[15][20] = 4'hE;
    SS5[16][20] = 4'hE;
    SS5[17][20] = 4'hE;
    SS5[18][20] = 4'hE;
    SS5[19][20] = 4'hD;
    SS5[20][20] = 4'hD;
    SS5[21][20] = 4'hD;
    SS5[22][20] = 4'hC;
    SS5[23][20] = 4'hC;
    SS5[24][20] = 4'hC;
    SS5[25][20] = 4'hC;
    SS5[26][20] = 4'hC;
    SS5[27][20] = 4'hC;
    SS5[28][20] = 4'hC;
    SS5[29][20] = 4'hD;
    SS5[30][20] = 4'hD;
    SS5[31][20] = 4'hD;
    SS5[32][20] = 4'h0;
    SS5[33][20] = 4'h0;
    SS5[34][20] = 4'h0;
    SS5[35][20] = 4'h0;
    SS5[36][20] = 4'h0;
    SS5[37][20] = 4'h0;
    SS5[38][20] = 4'h0;
    SS5[39][20] = 4'h0;
    SS5[40][20] = 4'h0;
    SS5[41][20] = 4'h0;
    SS5[42][20] = 4'h0;
    SS5[43][20] = 4'h0;
    SS5[44][20] = 4'h0;
    SS5[45][20] = 4'h0;
    SS5[46][20] = 4'h0;
    SS5[47][20] = 4'h0;
    SS5[0][21] = 4'h0;
    SS5[1][21] = 4'h0;
    SS5[2][21] = 4'h0;
    SS5[3][21] = 4'h0;
    SS5[4][21] = 4'h0;
    SS5[5][21] = 4'h0;
    SS5[6][21] = 4'h0;
    SS5[7][21] = 4'h0;
    SS5[8][21] = 4'h0;
    SS5[9][21] = 4'hE;
    SS5[10][21] = 4'h0;
    SS5[11][21] = 4'h0;
    SS5[12][21] = 4'hE;
    SS5[13][21] = 4'hE;
    SS5[14][21] = 4'hE;
    SS5[15][21] = 4'hE;
    SS5[16][21] = 4'hE;
    SS5[17][21] = 4'hE;
    SS5[18][21] = 4'hE;
    SS5[19][21] = 4'hD;
    SS5[20][21] = 4'hD;
    SS5[21][21] = 4'hD;
    SS5[22][21] = 4'hC;
    SS5[23][21] = 4'hC;
    SS5[24][21] = 4'hC;
    SS5[25][21] = 4'hD;
    SS5[26][21] = 4'hC;
    SS5[27][21] = 4'hC;
    SS5[28][21] = 4'hD;
    SS5[29][21] = 4'hD;
    SS5[30][21] = 4'hD;
    SS5[31][21] = 4'hC;
    SS5[32][21] = 4'hC;
    SS5[33][21] = 4'hE;
    SS5[34][21] = 4'h0;
    SS5[35][21] = 4'h0;
    SS5[36][21] = 4'h0;
    SS5[37][21] = 4'h0;
    SS5[38][21] = 4'h0;
    SS5[39][21] = 4'h0;
    SS5[40][21] = 4'h0;
    SS5[41][21] = 4'h0;
    SS5[42][21] = 4'h0;
    SS5[43][21] = 4'h0;
    SS5[44][21] = 4'h0;
    SS5[45][21] = 4'h0;
    SS5[46][21] = 4'h0;
    SS5[47][21] = 4'h0;
    SS5[0][22] = 4'h0;
    SS5[1][22] = 4'h0;
    SS5[2][22] = 4'h0;
    SS5[3][22] = 4'h0;
    SS5[4][22] = 4'h0;
    SS5[5][22] = 4'h0;
    SS5[6][22] = 4'h0;
    SS5[7][22] = 4'h0;
    SS5[8][22] = 4'h0;
    SS5[9][22] = 4'hE;
    SS5[10][22] = 4'hE;
    SS5[11][22] = 4'hE;
    SS5[12][22] = 4'hD;
    SS5[13][22] = 4'hE;
    SS5[14][22] = 4'hE;
    SS5[15][22] = 4'hE;
    SS5[16][22] = 4'hE;
    SS5[17][22] = 4'hE;
    SS5[18][22] = 4'hD;
    SS5[19][22] = 4'hD;
    SS5[20][22] = 4'hD;
    SS5[21][22] = 4'hC;
    SS5[22][22] = 4'hC;
    SS5[23][22] = 4'hC;
    SS5[24][22] = 4'hC;
    SS5[25][22] = 4'hD;
    SS5[26][22] = 4'hD;
    SS5[27][22] = 4'hD;
    SS5[28][22] = 4'hD;
    SS5[29][22] = 4'hD;
    SS5[30][22] = 4'hD;
    SS5[31][22] = 4'hC;
    SS5[32][22] = 4'hC;
    SS5[33][22] = 4'hC;
    SS5[34][22] = 4'hD;
    SS5[35][22] = 4'hD;
    SS5[36][22] = 4'h0;
    SS5[37][22] = 4'h0;
    SS5[38][22] = 4'h0;
    SS5[39][22] = 4'h0;
    SS5[40][22] = 4'h0;
    SS5[41][22] = 4'h0;
    SS5[42][22] = 4'h0;
    SS5[43][22] = 4'h0;
    SS5[44][22] = 4'h0;
    SS5[45][22] = 4'h0;
    SS5[46][22] = 4'h0;
    SS5[47][22] = 4'h0;
    SS5[0][23] = 4'h0;
    SS5[1][23] = 4'h0;
    SS5[2][23] = 4'h0;
    SS5[3][23] = 4'h0;
    SS5[4][23] = 4'h0;
    SS5[5][23] = 4'hE;
    SS5[6][23] = 4'hE;
    SS5[7][23] = 4'h0;
    SS5[8][23] = 4'hE;
    SS5[9][23] = 4'hE;
    SS5[10][23] = 4'hE;
    SS5[11][23] = 4'hD;
    SS5[12][23] = 4'hD;
    SS5[13][23] = 4'hD;
    SS5[14][23] = 4'hD;
    SS5[15][23] = 4'hE;
    SS5[16][23] = 4'hE;
    SS5[17][23] = 4'hE;
    SS5[18][23] = 4'hD;
    SS5[19][23] = 4'hD;
    SS5[20][23] = 4'hD;
    SS5[21][23] = 4'hC;
    SS5[22][23] = 4'hC;
    SS5[23][23] = 4'hC;
    SS5[24][23] = 4'hD;
    SS5[25][23] = 4'hD;
    SS5[26][23] = 4'hD;
    SS5[27][23] = 4'hA;
    SS5[28][23] = 4'hA;
    SS5[29][23] = 4'hA;
    SS5[30][23] = 4'hA;
    SS5[31][23] = 4'hC;
    SS5[32][23] = 4'hC;
    SS5[33][23] = 4'hC;
    SS5[34][23] = 4'hD;
    SS5[35][23] = 4'hD;
    SS5[36][23] = 4'hD;
    SS5[37][23] = 4'hD;
    SS5[38][23] = 4'h0;
    SS5[39][23] = 4'h0;
    SS5[40][23] = 4'h0;
    SS5[41][23] = 4'h0;
    SS5[42][23] = 4'h0;
    SS5[43][23] = 4'h0;
    SS5[44][23] = 4'h0;
    SS5[45][23] = 4'h0;
    SS5[46][23] = 4'h0;
    SS5[47][23] = 4'h0;
    SS5[0][24] = 4'h0;
    SS5[1][24] = 4'hD;
    SS5[2][24] = 4'h0;
    SS5[3][24] = 4'h0;
    SS5[4][24] = 4'h0;
    SS5[5][24] = 4'hE;
    SS5[6][24] = 4'hE;
    SS5[7][24] = 4'hE;
    SS5[8][24] = 4'hD;
    SS5[9][24] = 4'hD;
    SS5[10][24] = 4'hE;
    SS5[11][24] = 4'hD;
    SS5[12][24] = 4'hD;
    SS5[13][24] = 4'hD;
    SS5[14][24] = 4'hC;
    SS5[15][24] = 4'hC;
    SS5[16][24] = 4'hC;
    SS5[17][24] = 4'hD;
    SS5[18][24] = 4'hD;
    SS5[19][24] = 4'hD;
    SS5[20][24] = 4'hD;
    SS5[21][24] = 4'hC;
    SS5[22][24] = 4'hC;
    SS5[23][24] = 4'hC;
    SS5[24][24] = 4'hD;
    SS5[25][24] = 4'hD;
    SS5[26][24] = 4'hD;
    SS5[27][24] = 4'hA;
    SS5[28][24] = 4'hA;
    SS5[29][24] = 4'hA;
    SS5[30][24] = 4'hC;
    SS5[31][24] = 4'hC;
    SS5[32][24] = 4'hC;
    SS5[33][24] = 4'hD;
    SS5[34][24] = 4'hD;
    SS5[35][24] = 4'hD;
    SS5[36][24] = 4'hD;
    SS5[37][24] = 4'hD;
    SS5[38][24] = 4'hD;
    SS5[39][24] = 4'hD;
    SS5[40][24] = 4'hD;
    SS5[41][24] = 4'h0;
    SS5[42][24] = 4'h0;
    SS5[43][24] = 4'h0;
    SS5[44][24] = 4'h0;
    SS5[45][24] = 4'h0;
    SS5[46][24] = 4'h0;
    SS5[47][24] = 4'h0;
    SS5[0][25] = 4'h0;
    SS5[1][25] = 4'hD;
    SS5[2][25] = 4'hD;
    SS5[3][25] = 4'hD;
    SS5[4][25] = 4'hE;
    SS5[5][25] = 4'hE;
    SS5[6][25] = 4'hE;
    SS5[7][25] = 4'hD;
    SS5[8][25] = 4'hD;
    SS5[9][25] = 4'hD;
    SS5[10][25] = 4'hD;
    SS5[11][25] = 4'hC;
    SS5[12][25] = 4'hD;
    SS5[13][25] = 4'hD;
    SS5[14][25] = 4'hC;
    SS5[15][25] = 4'hC;
    SS5[16][25] = 4'hC;
    SS5[17][25] = 4'hC;
    SS5[18][25] = 4'hC;
    SS5[19][25] = 4'hC;
    SS5[20][25] = 4'hC;
    SS5[21][25] = 4'hC;
    SS5[22][25] = 4'hC;
    SS5[23][25] = 4'hD;
    SS5[24][25] = 4'hD;
    SS5[25][25] = 4'hD;
    SS5[26][25] = 4'hD;
    SS5[27][25] = 4'hA;
    SS5[28][25] = 4'hA;
    SS5[29][25] = 4'hA;
    SS5[30][25] = 4'hC;
    SS5[31][25] = 4'hC;
    SS5[32][25] = 4'hC;
    SS5[33][25] = 4'hC;
    SS5[34][25] = 4'hC;
    SS5[35][25] = 4'hD;
    SS5[36][25] = 4'hD;
    SS5[37][25] = 4'hD;
    SS5[38][25] = 4'hD;
    SS5[39][25] = 4'hD;
    SS5[40][25] = 4'hD;
    SS5[41][25] = 4'hD;
    SS5[42][25] = 4'hD;
    SS5[43][25] = 4'h0;
    SS5[44][25] = 4'h0;
    SS5[45][25] = 4'h0;
    SS5[46][25] = 4'h0;
    SS5[47][25] = 4'h0;
    SS5[0][26] = 4'h0;
    SS5[1][26] = 4'hD;
    SS5[2][26] = 4'hD;
    SS5[3][26] = 4'hD;
    SS5[4][26] = 4'hC;
    SS5[5][26] = 4'hC;
    SS5[6][26] = 4'hC;
    SS5[7][26] = 4'hD;
    SS5[8][26] = 4'hD;
    SS5[9][26] = 4'hD;
    SS5[10][26] = 4'hC;
    SS5[11][26] = 4'hC;
    SS5[12][26] = 4'hC;
    SS5[13][26] = 4'hC;
    SS5[14][26] = 4'hC;
    SS5[15][26] = 4'hC;
    SS5[16][26] = 4'hC;
    SS5[17][26] = 4'hC;
    SS5[18][26] = 4'hC;
    SS5[19][26] = 4'hC;
    SS5[20][26] = 4'hC;
    SS5[21][26] = 4'hC;
    SS5[22][26] = 4'hC;
    SS5[23][26] = 4'hD;
    SS5[24][26] = 4'hD;
    SS5[25][26] = 4'hD;
    SS5[26][26] = 4'hA;
    SS5[27][26] = 4'hA;
    SS5[28][26] = 4'hA;
    SS5[29][26] = 4'hC;
    SS5[30][26] = 4'hC;
    SS5[31][26] = 4'hC;
    SS5[32][26] = 4'hC;
    SS5[33][26] = 4'hC;
    SS5[34][26] = 4'hC;
    SS5[35][26] = 4'hC;
    SS5[36][26] = 4'hC;
    SS5[37][26] = 4'hC;
    SS5[38][26] = 4'hD;
    SS5[39][26] = 4'hD;
    SS5[40][26] = 4'hD;
    SS5[41][26] = 4'hD;
    SS5[42][26] = 4'h0;
    SS5[43][26] = 4'h0;
    SS5[44][26] = 4'h0;
    SS5[45][26] = 4'h0;
    SS5[46][26] = 4'h0;
    SS5[47][26] = 4'h0;
    SS5[0][27] = 4'hC;
    SS5[1][27] = 4'hD;
    SS5[2][27] = 4'hD;
    SS5[3][27] = 4'hC;
    SS5[4][27] = 4'hC;
    SS5[5][27] = 4'hC;
    SS5[6][27] = 4'hC;
    SS5[7][27] = 4'hC;
    SS5[8][27] = 4'hC;
    SS5[9][27] = 4'hD;
    SS5[10][27] = 4'hC;
    SS5[11][27] = 4'hC;
    SS5[12][27] = 4'hC;
    SS5[13][27] = 4'hC;
    SS5[14][27] = 4'hC;
    SS5[15][27] = 4'hC;
    SS5[16][27] = 4'hC;
    SS5[17][27] = 4'hC;
    SS5[18][27] = 4'hC;
    SS5[19][27] = 4'hC;
    SS5[20][27] = 4'hC;
    SS5[21][27] = 4'hC;
    SS5[22][27] = 4'hC;
    SS5[23][27] = 4'hC;
    SS5[24][27] = 4'hC;
    SS5[25][27] = 4'hD;
    SS5[26][27] = 4'hA;
    SS5[27][27] = 4'hA;
    SS5[28][27] = 4'hA;
    SS5[29][27] = 4'hC;
    SS5[30][27] = 4'hC;
    SS5[31][27] = 4'hC;
    SS5[32][27] = 4'hC;
    SS5[33][27] = 4'hC;
    SS5[34][27] = 4'hC;
    SS5[35][27] = 4'hC;
    SS5[36][27] = 4'hC;
    SS5[37][27] = 4'hC;
    SS5[38][27] = 4'hC;
    SS5[39][27] = 4'hC;
    SS5[40][27] = 4'hD;
    SS5[41][27] = 4'hD;
    SS5[42][27] = 4'h0;
    SS5[43][27] = 4'h0;
    SS5[44][27] = 4'h0;
    SS5[45][27] = 4'h0;
    SS5[46][27] = 4'h0;
    SS5[47][27] = 4'h0;
    SS5[0][28] = 4'hC;
    SS5[1][28] = 4'hC;
    SS5[2][28] = 4'hC;
    SS5[3][28] = 4'hC;
    SS5[4][28] = 4'hC;
    SS5[5][28] = 4'hC;
    SS5[6][28] = 4'hC;
    SS5[7][28] = 4'hC;
    SS5[8][28] = 4'hC;
    SS5[9][28] = 4'hC;
    SS5[10][28] = 4'hC;
    SS5[11][28] = 4'hC;
    SS5[12][28] = 4'hC;
    SS5[13][28] = 4'hC;
    SS5[14][28] = 4'hC;
    SS5[15][28] = 4'hC;
    SS5[16][28] = 4'hC;
    SS5[17][28] = 4'hC;
    SS5[18][28] = 4'hC;
    SS5[19][28] = 4'hC;
    SS5[20][28] = 4'hC;
    SS5[21][28] = 4'hC;
    SS5[22][28] = 4'hC;
    SS5[23][28] = 4'hC;
    SS5[24][28] = 4'hC;
    SS5[25][28] = 4'hD;
    SS5[26][28] = 4'hD;
    SS5[27][28] = 4'hA;
    SS5[28][28] = 4'hA;
    SS5[29][28] = 4'hC;
    SS5[30][28] = 4'hC;
    SS5[31][28] = 4'hC;
    SS5[32][28] = 4'hC;
    SS5[33][28] = 4'hC;
    SS5[34][28] = 4'hC;
    SS5[35][28] = 4'hC;
    SS5[36][28] = 4'hC;
    SS5[37][28] = 4'hC;
    SS5[38][28] = 4'hC;
    SS5[39][28] = 4'hC;
    SS5[40][28] = 4'hC;
    SS5[41][28] = 4'hC;
    SS5[42][28] = 4'hC;
    SS5[43][28] = 4'h0;
    SS5[44][28] = 4'h0;
    SS5[45][28] = 4'h0;
    SS5[46][28] = 4'h0;
    SS5[47][28] = 4'h0;
    SS5[0][29] = 4'hC;
    SS5[1][29] = 4'hC;
    SS5[2][29] = 4'hC;
    SS5[3][29] = 4'hC;
    SS5[4][29] = 4'hC;
    SS5[5][29] = 4'hC;
    SS5[6][29] = 4'hC;
    SS5[7][29] = 4'hC;
    SS5[8][29] = 4'hC;
    SS5[9][29] = 4'hC;
    SS5[10][29] = 4'hC;
    SS5[11][29] = 4'hC;
    SS5[12][29] = 4'hC;
    SS5[13][29] = 4'hC;
    SS5[14][29] = 4'hC;
    SS5[15][29] = 4'hC;
    SS5[16][29] = 4'hC;
    SS5[17][29] = 4'hC;
    SS5[18][29] = 4'hC;
    SS5[19][29] = 4'hE;
    SS5[20][29] = 4'hE;
    SS5[21][29] = 4'hE;
    SS5[22][29] = 4'hC;
    SS5[23][29] = 4'hC;
    SS5[24][29] = 4'hC;
    SS5[25][29] = 4'hD;
    SS5[26][29] = 4'hD;
    SS5[27][29] = 4'hD;
    SS5[28][29] = 4'hC;
    SS5[29][29] = 4'hC;
    SS5[30][29] = 4'hC;
    SS5[31][29] = 4'hC;
    SS5[32][29] = 4'hC;
    SS5[33][29] = 4'hC;
    SS5[34][29] = 4'hC;
    SS5[35][29] = 4'hC;
    SS5[36][29] = 4'hC;
    SS5[37][29] = 4'hC;
    SS5[38][29] = 4'hC;
    SS5[39][29] = 4'hC;
    SS5[40][29] = 4'hC;
    SS5[41][29] = 4'hC;
    SS5[42][29] = 4'hC;
    SS5[43][29] = 4'hC;
    SS5[44][29] = 4'hC;
    SS5[45][29] = 4'h0;
    SS5[46][29] = 4'h0;
    SS5[47][29] = 4'h0;
    SS5[0][30] = 4'h0;
    SS5[1][30] = 4'hC;
    SS5[2][30] = 4'hC;
    SS5[3][30] = 4'hC;
    SS5[4][30] = 4'hC;
    SS5[5][30] = 4'h0;
    SS5[6][30] = 4'h0;
    SS5[7][30] = 4'h0;
    SS5[8][30] = 4'h0;
    SS5[9][30] = 4'hC;
    SS5[10][30] = 4'hC;
    SS5[11][30] = 4'hC;
    SS5[12][30] = 4'hC;
    SS5[13][30] = 4'hC;
    SS5[14][30] = 4'hC;
    SS5[15][30] = 4'hE;
    SS5[16][30] = 4'hC;
    SS5[17][30] = 4'hC;
    SS5[18][30] = 4'hE;
    SS5[19][30] = 4'hE;
    SS5[20][30] = 4'hE;
    SS5[21][30] = 4'hD;
    SS5[22][30] = 4'hD;
    SS5[23][30] = 4'hD;
    SS5[24][30] = 4'hC;
    SS5[25][30] = 4'hD;
    SS5[26][30] = 4'hD;
    SS5[27][30] = 4'hD;
    SS5[28][30] = 4'hC;
    SS5[29][30] = 4'hC;
    SS5[30][30] = 4'hC;
    SS5[31][30] = 4'hD;
    SS5[32][30] = 4'hC;
    SS5[33][30] = 4'hC;
    SS5[34][30] = 4'hC;
    SS5[35][30] = 4'hC;
    SS5[36][30] = 4'hC;
    SS5[37][30] = 4'hC;
    SS5[38][30] = 4'hC;
    SS5[39][30] = 4'hC;
    SS5[40][30] = 4'hC;
    SS5[41][30] = 4'hC;
    SS5[42][30] = 4'hC;
    SS5[43][30] = 4'hC;
    SS5[44][30] = 4'hC;
    SS5[45][30] = 4'hC;
    SS5[46][30] = 4'hC;
    SS5[47][30] = 4'h0;
    SS5[0][31] = 4'h0;
    SS5[1][31] = 4'h0;
    SS5[2][31] = 4'h0;
    SS5[3][31] = 4'hC;
    SS5[4][31] = 4'hC;
    SS5[5][31] = 4'h0;
    SS5[6][31] = 4'h0;
    SS5[7][31] = 4'h0;
    SS5[8][31] = 4'h0;
    SS5[9][31] = 4'h0;
    SS5[10][31] = 4'h0;
    SS5[11][31] = 4'hC;
    SS5[12][31] = 4'hC;
    SS5[13][31] = 4'hC;
    SS5[14][31] = 4'hE;
    SS5[15][31] = 4'hE;
    SS5[16][31] = 4'hE;
    SS5[17][31] = 4'hE;
    SS5[18][31] = 4'hD;
    SS5[19][31] = 4'hE;
    SS5[20][31] = 4'hE;
    SS5[21][31] = 4'hD;
    SS5[22][31] = 4'hD;
    SS5[23][31] = 4'hD;
    SS5[24][31] = 4'hD;
    SS5[25][31] = 4'hD;
    SS5[26][31] = 4'hD;
    SS5[27][31] = 4'hC;
    SS5[28][31] = 4'hC;
    SS5[29][31] = 4'hC;
    SS5[30][31] = 4'hC;
    SS5[31][31] = 4'hD;
    SS5[32][31] = 4'hD;
    SS5[33][31] = 4'hD;
    SS5[34][31] = 4'hC;
    SS5[35][31] = 4'hC;
    SS5[36][31] = 4'hC;
    SS5[37][31] = 4'hC;
    SS5[38][31] = 4'hC;
    SS5[39][31] = 4'hC;
    SS5[40][31] = 4'hC;
    SS5[41][31] = 4'hC;
    SS5[42][31] = 4'hC;
    SS5[43][31] = 4'hC;
    SS5[44][31] = 4'hC;
    SS5[45][31] = 4'hC;
    SS5[46][31] = 4'hC;
    SS5[47][31] = 4'h0;
    SS5[0][32] = 4'h0;
    SS5[1][32] = 4'h0;
    SS5[2][32] = 4'h0;
    SS5[3][32] = 4'h0;
    SS5[4][32] = 4'h0;
    SS5[5][32] = 4'h0;
    SS5[6][32] = 4'h0;
    SS5[7][32] = 4'h0;
    SS5[8][32] = 4'h0;
    SS5[9][32] = 4'h0;
    SS5[10][32] = 4'h0;
    SS5[11][32] = 4'hE;
    SS5[12][32] = 4'hE;
    SS5[13][32] = 4'hE;
    SS5[14][32] = 4'hE;
    SS5[15][32] = 4'hE;
    SS5[16][32] = 4'hE;
    SS5[17][32] = 4'hD;
    SS5[18][32] = 4'hD;
    SS5[19][32] = 4'hD;
    SS5[20][32] = 4'hD;
    SS5[21][32] = 4'hD;
    SS5[22][32] = 4'hD;
    SS5[23][32] = 4'hD;
    SS5[24][32] = 4'hD;
    SS5[25][32] = 4'hD;
    SS5[26][32] = 4'hD;
    SS5[27][32] = 4'h0;
    SS5[28][32] = 4'h0;
    SS5[29][32] = 4'hC;
    SS5[30][32] = 4'hD;
    SS5[31][32] = 4'hD;
    SS5[32][32] = 4'hD;
    SS5[33][32] = 4'hD;
    SS5[34][32] = 4'hD;
    SS5[35][32] = 4'hD;
    SS5[36][32] = 4'hD;
    SS5[37][32] = 4'hC;
    SS5[38][32] = 4'hC;
    SS5[39][32] = 4'hC;
    SS5[40][32] = 4'hC;
    SS5[41][32] = 4'hC;
    SS5[42][32] = 4'hC;
    SS5[43][32] = 4'hC;
    SS5[44][32] = 4'hC;
    SS5[45][32] = 4'hC;
    SS5[46][32] = 4'h0;
    SS5[47][32] = 4'h0;
    SS5[0][33] = 4'h0;
    SS5[1][33] = 4'h0;
    SS5[2][33] = 4'h0;
    SS5[3][33] = 4'h0;
    SS5[4][33] = 4'h0;
    SS5[5][33] = 4'h0;
    SS5[6][33] = 4'h0;
    SS5[7][33] = 4'h0;
    SS5[8][33] = 4'h0;
    SS5[9][33] = 4'h0;
    SS5[10][33] = 4'hE;
    SS5[11][33] = 4'hE;
    SS5[12][33] = 4'hE;
    SS5[13][33] = 4'hE;
    SS5[14][33] = 4'hE;
    SS5[15][33] = 4'hE;
    SS5[16][33] = 4'hE;
    SS5[17][33] = 4'hD;
    SS5[18][33] = 4'hD;
    SS5[19][33] = 4'hD;
    SS5[20][33] = 4'hD;
    SS5[21][33] = 4'hD;
    SS5[22][33] = 4'hD;
    SS5[23][33] = 4'h3;
    SS5[24][33] = 4'hD;
    SS5[25][33] = 4'hD;
    SS5[26][33] = 4'hF;
    SS5[27][33] = 4'h0;
    SS5[28][33] = 4'h0;
    SS5[29][33] = 4'h0;
    SS5[30][33] = 4'h0;
    SS5[31][33] = 4'hD;
    SS5[32][33] = 4'hD;
    SS5[33][33] = 4'hD;
    SS5[34][33] = 4'hD;
    SS5[35][33] = 4'hD;
    SS5[36][33] = 4'hD;
    SS5[37][33] = 4'hD;
    SS5[38][33] = 4'hD;
    SS5[39][33] = 4'hC;
    SS5[40][33] = 4'hC;
    SS5[41][33] = 4'hC;
    SS5[42][33] = 4'hC;
    SS5[43][33] = 4'hC;
    SS5[44][33] = 4'hC;
    SS5[45][33] = 4'hC;
    SS5[46][33] = 4'h0;
    SS5[47][33] = 4'h0;
    SS5[0][34] = 4'h0;
    SS5[1][34] = 4'h0;
    SS5[2][34] = 4'h0;
    SS5[3][34] = 4'h0;
    SS5[4][34] = 4'h0;
    SS5[5][34] = 4'h0;
    SS5[6][34] = 4'h0;
    SS5[7][34] = 4'h0;
    SS5[8][34] = 4'h0;
    SS5[9][34] = 4'h0;
    SS5[10][34] = 4'hE;
    SS5[11][34] = 4'hE;
    SS5[12][34] = 4'hE;
    SS5[13][34] = 4'hE;
    SS5[14][34] = 4'hE;
    SS5[15][34] = 4'hE;
    SS5[16][34] = 4'hD;
    SS5[17][34] = 4'hD;
    SS5[18][34] = 4'hD;
    SS5[19][34] = 4'hD;
    SS5[20][34] = 4'hD;
    SS5[21][34] = 4'hD;
    SS5[22][34] = 4'hD;
    SS5[23][34] = 4'h3;
    SS5[24][34] = 4'h3;
    SS5[25][34] = 4'h3;
    SS5[26][34] = 4'h0;
    SS5[27][34] = 4'h0;
    SS5[28][34] = 4'h0;
    SS5[29][34] = 4'h0;
    SS5[30][34] = 4'h0;
    SS5[31][34] = 4'h0;
    SS5[32][34] = 4'h0;
    SS5[33][34] = 4'h0;
    SS5[34][34] = 4'hD;
    SS5[35][34] = 4'hD;
    SS5[36][34] = 4'hD;
    SS5[37][34] = 4'hD;
    SS5[38][34] = 4'hD;
    SS5[39][34] = 4'h0;
    SS5[40][34] = 4'h0;
    SS5[41][34] = 4'h0;
    SS5[42][34] = 4'hC;
    SS5[43][34] = 4'hC;
    SS5[44][34] = 4'hC;
    SS5[45][34] = 4'h0;
    SS5[46][34] = 4'h0;
    SS5[47][34] = 4'h0;
    SS5[0][35] = 4'h0;
    SS5[1][35] = 4'h0;
    SS5[2][35] = 4'h0;
    SS5[3][35] = 4'h0;
    SS5[4][35] = 4'h0;
    SS5[5][35] = 4'h0;
    SS5[6][35] = 4'h0;
    SS5[7][35] = 4'h0;
    SS5[8][35] = 4'h0;
    SS5[9][35] = 4'h0;
    SS5[10][35] = 4'hE;
    SS5[11][35] = 4'hE;
    SS5[12][35] = 4'hE;
    SS5[13][35] = 4'hE;
    SS5[14][35] = 4'hE;
    SS5[15][35] = 4'hE;
    SS5[16][35] = 4'hD;
    SS5[17][35] = 4'hD;
    SS5[18][35] = 4'hD;
    SS5[19][35] = 4'h0;
    SS5[20][35] = 4'h0;
    SS5[21][35] = 4'hD;
    SS5[22][35] = 4'h3;
    SS5[23][35] = 4'h3;
    SS5[24][35] = 4'h3;
    SS5[25][35] = 4'h3;
    SS5[26][35] = 4'h0;
    SS5[27][35] = 4'h0;
    SS5[28][35] = 4'h0;
    SS5[29][35] = 4'h0;
    SS5[30][35] = 4'h0;
    SS5[31][35] = 4'h0;
    SS5[32][35] = 4'h0;
    SS5[33][35] = 4'h0;
    SS5[34][35] = 4'h0;
    SS5[35][35] = 4'h0;
    SS5[36][35] = 4'hD;
    SS5[37][35] = 4'hD;
    SS5[38][35] = 4'hF;
    SS5[39][35] = 4'h0;
    SS5[40][35] = 4'h0;
    SS5[41][35] = 4'h0;
    SS5[42][35] = 4'h0;
    SS5[43][35] = 4'h0;
    SS5[44][35] = 4'hC;
    SS5[45][35] = 4'h0;
    SS5[46][35] = 4'h0;
    SS5[47][35] = 4'h0;
    SS5[0][36] = 4'h0;
    SS5[1][36] = 4'h0;
    SS5[2][36] = 4'h0;
    SS5[3][36] = 4'h0;
    SS5[4][36] = 4'h0;
    SS5[5][36] = 4'h0;
    SS5[6][36] = 4'h0;
    SS5[7][36] = 4'h0;
    SS5[8][36] = 4'h0;
    SS5[9][36] = 4'hE;
    SS5[10][36] = 4'hE;
    SS5[11][36] = 4'hE;
    SS5[12][36] = 4'hD;
    SS5[13][36] = 4'hD;
    SS5[14][36] = 4'hD;
    SS5[15][36] = 4'hE;
    SS5[16][36] = 4'hD;
    SS5[17][36] = 4'hD;
    SS5[18][36] = 4'hD;
    SS5[19][36] = 4'h0;
    SS5[20][36] = 4'h0;
    SS5[21][36] = 4'h0;
    SS5[22][36] = 4'h0;
    SS5[23][36] = 4'h3;
    SS5[24][36] = 4'h3;
    SS5[25][36] = 4'h0;
    SS5[26][36] = 4'h0;
    SS5[27][36] = 4'h0;
    SS5[28][36] = 4'h0;
    SS5[29][36] = 4'h0;
    SS5[30][36] = 4'h0;
    SS5[31][36] = 4'h0;
    SS5[32][36] = 4'h0;
    SS5[33][36] = 4'h0;
    SS5[34][36] = 4'h0;
    SS5[35][36] = 4'h0;
    SS5[36][36] = 4'h0;
    SS5[37][36] = 4'h0;
    SS5[38][36] = 4'h0;
    SS5[39][36] = 4'h0;
    SS5[40][36] = 4'h0;
    SS5[41][36] = 4'h0;
    SS5[42][36] = 4'h0;
    SS5[43][36] = 4'h0;
    SS5[44][36] = 4'h0;
    SS5[45][36] = 4'h0;
    SS5[46][36] = 4'h0;
    SS5[47][36] = 4'h0;
    SS5[0][37] = 4'h0;
    SS5[1][37] = 4'h0;
    SS5[2][37] = 4'h0;
    SS5[3][37] = 4'h0;
    SS5[4][37] = 4'h0;
    SS5[5][37] = 4'h0;
    SS5[6][37] = 4'h0;
    SS5[7][37] = 4'h0;
    SS5[8][37] = 4'h0;
    SS5[9][37] = 4'hD;
    SS5[10][37] = 4'hE;
    SS5[11][37] = 4'hE;
    SS5[12][37] = 4'hD;
    SS5[13][37] = 4'hD;
    SS5[14][37] = 4'hD;
    SS5[15][37] = 4'h3;
    SS5[16][37] = 4'h3;
    SS5[17][37] = 4'h3;
    SS5[18][37] = 4'h0;
    SS5[19][37] = 4'h0;
    SS5[20][37] = 4'h0;
    SS5[21][37] = 4'h0;
    SS5[22][37] = 4'h0;
    SS5[23][37] = 4'h0;
    SS5[24][37] = 4'h0;
    SS5[25][37] = 4'h0;
    SS5[26][37] = 4'h0;
    SS5[27][37] = 4'h0;
    SS5[28][37] = 4'h0;
    SS5[29][37] = 4'h0;
    SS5[30][37] = 4'h0;
    SS5[31][37] = 4'h0;
    SS5[32][37] = 4'h0;
    SS5[33][37] = 4'h0;
    SS5[34][37] = 4'h0;
    SS5[35][37] = 4'h0;
    SS5[36][37] = 4'h0;
    SS5[37][37] = 4'h0;
    SS5[38][37] = 4'h0;
    SS5[39][37] = 4'h0;
    SS5[40][37] = 4'h0;
    SS5[41][37] = 4'h0;
    SS5[42][37] = 4'h0;
    SS5[43][37] = 4'h0;
    SS5[44][37] = 4'h0;
    SS5[45][37] = 4'h0;
    SS5[46][37] = 4'h0;
    SS5[47][37] = 4'h0;
    SS5[0][38] = 4'h0;
    SS5[1][38] = 4'h0;
    SS5[2][38] = 4'h0;
    SS5[3][38] = 4'h0;
    SS5[4][38] = 4'h0;
    SS5[5][38] = 4'h0;
    SS5[6][38] = 4'h0;
    SS5[7][38] = 4'h0;
    SS5[8][38] = 4'hD;
    SS5[9][38] = 4'hD;
    SS5[10][38] = 4'hD;
    SS5[11][38] = 4'hD;
    SS5[12][38] = 4'hD;
    SS5[13][38] = 4'hD;
    SS5[14][38] = 4'hD;
    SS5[15][38] = 4'h3;
    SS5[16][38] = 4'h3;
    SS5[17][38] = 4'h3;
    SS5[18][38] = 4'h0;
    SS5[19][38] = 4'h0;
    SS5[20][38] = 4'h0;
    SS5[21][38] = 4'h0;
    SS5[22][38] = 4'h0;
    SS5[23][38] = 4'h0;
    SS5[24][38] = 4'h0;
    SS5[25][38] = 4'h0;
    SS5[26][38] = 4'h0;
    SS5[27][38] = 4'h0;
    SS5[28][38] = 4'h0;
    SS5[29][38] = 4'h0;
    SS5[30][38] = 4'h0;
    SS5[31][38] = 4'h0;
    SS5[32][38] = 4'h0;
    SS5[33][38] = 4'h0;
    SS5[34][38] = 4'h0;
    SS5[35][38] = 4'h0;
    SS5[36][38] = 4'h0;
    SS5[37][38] = 4'h0;
    SS5[38][38] = 4'h0;
    SS5[39][38] = 4'h0;
    SS5[40][38] = 4'h0;
    SS5[41][38] = 4'h0;
    SS5[42][38] = 4'h0;
    SS5[43][38] = 4'h0;
    SS5[44][38] = 4'h0;
    SS5[45][38] = 4'h0;
    SS5[46][38] = 4'h0;
    SS5[47][38] = 4'h0;
    SS5[0][39] = 4'h0;
    SS5[1][39] = 4'h0;
    SS5[2][39] = 4'h0;
    SS5[3][39] = 4'h0;
    SS5[4][39] = 4'h0;
    SS5[5][39] = 4'h0;
    SS5[6][39] = 4'h0;
    SS5[7][39] = 4'h0;
    SS5[8][39] = 4'hD;
    SS5[9][39] = 4'hD;
    SS5[10][39] = 4'hD;
    SS5[11][39] = 4'hD;
    SS5[12][39] = 4'hD;
    SS5[13][39] = 4'hD;
    SS5[14][39] = 4'h0;
    SS5[15][39] = 4'h3;
    SS5[16][39] = 4'h3;
    SS5[17][39] = 4'h3;
    SS5[18][39] = 4'h0;
    SS5[19][39] = 4'h0;
    SS5[20][39] = 4'h0;
    SS5[21][39] = 4'h0;
    SS5[22][39] = 4'h0;
    SS5[23][39] = 4'h0;
    SS5[24][39] = 4'h0;
    SS5[25][39] = 4'h0;
    SS5[26][39] = 4'h0;
    SS5[27][39] = 4'h0;
    SS5[28][39] = 4'h0;
    SS5[29][39] = 4'h0;
    SS5[30][39] = 4'h0;
    SS5[31][39] = 4'h0;
    SS5[32][39] = 4'h0;
    SS5[33][39] = 4'h0;
    SS5[34][39] = 4'h0;
    SS5[35][39] = 4'h0;
    SS5[36][39] = 4'h0;
    SS5[37][39] = 4'h0;
    SS5[38][39] = 4'h0;
    SS5[39][39] = 4'h0;
    SS5[40][39] = 4'h0;
    SS5[41][39] = 4'h0;
    SS5[42][39] = 4'h0;
    SS5[43][39] = 4'h0;
    SS5[44][39] = 4'h0;
    SS5[45][39] = 4'h0;
    SS5[46][39] = 4'h0;
    SS5[47][39] = 4'h0;
    SS5[0][40] = 4'h0;
    SS5[1][40] = 4'h0;
    SS5[2][40] = 4'h0;
    SS5[3][40] = 4'h0;
    SS5[4][40] = 4'h0;
    SS5[5][40] = 4'h0;
    SS5[6][40] = 4'h0;
    SS5[7][40] = 4'h0;
    SS5[8][40] = 4'hD;
    SS5[9][40] = 4'hD;
    SS5[10][40] = 4'hD;
    SS5[11][40] = 4'hD;
    SS5[12][40] = 4'hD;
    SS5[13][40] = 4'hD;
    SS5[14][40] = 4'h0;
    SS5[15][40] = 4'h0;
    SS5[16][40] = 4'h0;
    SS5[17][40] = 4'h0;
    SS5[18][40] = 4'h0;
    SS5[19][40] = 4'h0;
    SS5[20][40] = 4'h0;
    SS5[21][40] = 4'h0;
    SS5[22][40] = 4'h0;
    SS5[23][40] = 4'h0;
    SS5[24][40] = 4'h0;
    SS5[25][40] = 4'h0;
    SS5[26][40] = 4'h0;
    SS5[27][40] = 4'h0;
    SS5[28][40] = 4'h0;
    SS5[29][40] = 4'h0;
    SS5[30][40] = 4'h0;
    SS5[31][40] = 4'h0;
    SS5[32][40] = 4'h0;
    SS5[33][40] = 4'h0;
    SS5[34][40] = 4'h0;
    SS5[35][40] = 4'h0;
    SS5[36][40] = 4'h0;
    SS5[37][40] = 4'h0;
    SS5[38][40] = 4'h0;
    SS5[39][40] = 4'h0;
    SS5[40][40] = 4'h0;
    SS5[41][40] = 4'h0;
    SS5[42][40] = 4'h0;
    SS5[43][40] = 4'h0;
    SS5[44][40] = 4'h0;
    SS5[45][40] = 4'h0;
    SS5[46][40] = 4'h0;
    SS5[47][40] = 4'h0;
    SS5[0][41] = 4'h0;
    SS5[1][41] = 4'h0;
    SS5[2][41] = 4'h0;
    SS5[3][41] = 4'h0;
    SS5[4][41] = 4'h0;
    SS5[5][41] = 4'h0;
    SS5[6][41] = 4'h0;
    SS5[7][41] = 4'hD;
    SS5[8][41] = 4'hD;
    SS5[9][41] = 4'hD;
    SS5[10][41] = 4'h0;
    SS5[11][41] = 4'h0;
    SS5[12][41] = 4'hD;
    SS5[13][41] = 4'hD;
    SS5[14][41] = 4'h0;
    SS5[15][41] = 4'h0;
    SS5[16][41] = 4'h0;
    SS5[17][41] = 4'h0;
    SS5[18][41] = 4'h0;
    SS5[19][41] = 4'h0;
    SS5[20][41] = 4'h0;
    SS5[21][41] = 4'h0;
    SS5[22][41] = 4'h0;
    SS5[23][41] = 4'h0;
    SS5[24][41] = 4'h0;
    SS5[25][41] = 4'h0;
    SS5[26][41] = 4'h0;
    SS5[27][41] = 4'h0;
    SS5[28][41] = 4'h0;
    SS5[29][41] = 4'h0;
    SS5[30][41] = 4'h0;
    SS5[31][41] = 4'h0;
    SS5[32][41] = 4'h0;
    SS5[33][41] = 4'h0;
    SS5[34][41] = 4'h0;
    SS5[35][41] = 4'h0;
    SS5[36][41] = 4'h0;
    SS5[37][41] = 4'h0;
    SS5[38][41] = 4'h0;
    SS5[39][41] = 4'h0;
    SS5[40][41] = 4'h0;
    SS5[41][41] = 4'h0;
    SS5[42][41] = 4'h0;
    SS5[43][41] = 4'h0;
    SS5[44][41] = 4'h0;
    SS5[45][41] = 4'h0;
    SS5[46][41] = 4'h0;
    SS5[47][41] = 4'h0;
    SS5[0][42] = 4'h0;
    SS5[1][42] = 4'h0;
    SS5[2][42] = 4'h0;
    SS5[3][42] = 4'h0;
    SS5[4][42] = 4'h0;
    SS5[5][42] = 4'h0;
    SS5[6][42] = 4'h0;
    SS5[7][42] = 4'hD;
    SS5[8][42] = 4'hD;
    SS5[9][42] = 4'hD;
    SS5[10][42] = 4'h0;
    SS5[11][42] = 4'h0;
    SS5[12][42] = 4'h0;
    SS5[13][42] = 4'h0;
    SS5[14][42] = 4'h0;
    SS5[15][42] = 4'h0;
    SS5[16][42] = 4'h0;
    SS5[17][42] = 4'h0;
    SS5[18][42] = 4'h0;
    SS5[19][42] = 4'h0;
    SS5[20][42] = 4'h0;
    SS5[21][42] = 4'h0;
    SS5[22][42] = 4'h0;
    SS5[23][42] = 4'h0;
    SS5[24][42] = 4'h0;
    SS5[25][42] = 4'h0;
    SS5[26][42] = 4'h0;
    SS5[27][42] = 4'h0;
    SS5[28][42] = 4'h0;
    SS5[29][42] = 4'h0;
    SS5[30][42] = 4'h0;
    SS5[31][42] = 4'h0;
    SS5[32][42] = 4'h0;
    SS5[33][42] = 4'h0;
    SS5[34][42] = 4'h0;
    SS5[35][42] = 4'h0;
    SS5[36][42] = 4'h0;
    SS5[37][42] = 4'h0;
    SS5[38][42] = 4'h0;
    SS5[39][42] = 4'h0;
    SS5[40][42] = 4'h0;
    SS5[41][42] = 4'h0;
    SS5[42][42] = 4'h0;
    SS5[43][42] = 4'h0;
    SS5[44][42] = 4'h0;
    SS5[45][42] = 4'h0;
    SS5[46][42] = 4'h0;
    SS5[47][42] = 4'h0;
    SS5[0][43] = 4'h0;
    SS5[1][43] = 4'h0;
    SS5[2][43] = 4'h0;
    SS5[3][43] = 4'h0;
    SS5[4][43] = 4'h0;
    SS5[5][43] = 4'h0;
    SS5[6][43] = 4'h0;
    SS5[7][43] = 4'h0;
    SS5[8][43] = 4'h0;
    SS5[9][43] = 4'hD;
    SS5[10][43] = 4'h0;
    SS5[11][43] = 4'h0;
    SS5[12][43] = 4'h0;
    SS5[13][43] = 4'h0;
    SS5[14][43] = 4'h0;
    SS5[15][43] = 4'h0;
    SS5[16][43] = 4'h0;
    SS5[17][43] = 4'h0;
    SS5[18][43] = 4'h0;
    SS5[19][43] = 4'h0;
    SS5[20][43] = 4'h0;
    SS5[21][43] = 4'h0;
    SS5[22][43] = 4'h0;
    SS5[23][43] = 4'h0;
    SS5[24][43] = 4'h0;
    SS5[25][43] = 4'h0;
    SS5[26][43] = 4'h0;
    SS5[27][43] = 4'h0;
    SS5[28][43] = 4'h0;
    SS5[29][43] = 4'h0;
    SS5[30][43] = 4'h0;
    SS5[31][43] = 4'h0;
    SS5[32][43] = 4'h0;
    SS5[33][43] = 4'h0;
    SS5[34][43] = 4'h0;
    SS5[35][43] = 4'h0;
    SS5[36][43] = 4'h0;
    SS5[37][43] = 4'h0;
    SS5[38][43] = 4'h0;
    SS5[39][43] = 4'h0;
    SS5[40][43] = 4'h0;
    SS5[41][43] = 4'h0;
    SS5[42][43] = 4'h0;
    SS5[43][43] = 4'h0;
    SS5[44][43] = 4'h0;
    SS5[45][43] = 4'h0;
    SS5[46][43] = 4'h0;
    SS5[47][43] = 4'h0;
    SS5[0][44] = 4'h0;
    SS5[1][44] = 4'h0;
    SS5[2][44] = 4'h0;
    SS5[3][44] = 4'h0;
    SS5[4][44] = 4'h0;
    SS5[5][44] = 4'h0;
    SS5[6][44] = 4'h0;
    SS5[7][44] = 4'h0;
    SS5[8][44] = 4'h0;
    SS5[9][44] = 4'h0;
    SS5[10][44] = 4'h0;
    SS5[11][44] = 4'h0;
    SS5[12][44] = 4'h0;
    SS5[13][44] = 4'h0;
    SS5[14][44] = 4'h0;
    SS5[15][44] = 4'h0;
    SS5[16][44] = 4'h0;
    SS5[17][44] = 4'h0;
    SS5[18][44] = 4'h0;
    SS5[19][44] = 4'h0;
    SS5[20][44] = 4'h0;
    SS5[21][44] = 4'h0;
    SS5[22][44] = 4'h0;
    SS5[23][44] = 4'h0;
    SS5[24][44] = 4'h0;
    SS5[25][44] = 4'h0;
    SS5[26][44] = 4'h0;
    SS5[27][44] = 4'h0;
    SS5[28][44] = 4'h0;
    SS5[29][44] = 4'h0;
    SS5[30][44] = 4'h0;
    SS5[31][44] = 4'h0;
    SS5[32][44] = 4'h0;
    SS5[33][44] = 4'h0;
    SS5[34][44] = 4'h0;
    SS5[35][44] = 4'h0;
    SS5[36][44] = 4'h0;
    SS5[37][44] = 4'h0;
    SS5[38][44] = 4'h0;
    SS5[39][44] = 4'h0;
    SS5[40][44] = 4'h0;
    SS5[41][44] = 4'h0;
    SS5[42][44] = 4'h0;
    SS5[43][44] = 4'h0;
    SS5[44][44] = 4'h0;
    SS5[45][44] = 4'h0;
    SS5[46][44] = 4'h0;
    SS5[47][44] = 4'h0;
    SS5[0][45] = 4'h0;
    SS5[1][45] = 4'h0;
    SS5[2][45] = 4'h0;
    SS5[3][45] = 4'h0;
    SS5[4][45] = 4'h0;
    SS5[5][45] = 4'h0;
    SS5[6][45] = 4'h0;
    SS5[7][45] = 4'h0;
    SS5[8][45] = 4'h0;
    SS5[9][45] = 4'h0;
    SS5[10][45] = 4'h0;
    SS5[11][45] = 4'h0;
    SS5[12][45] = 4'h0;
    SS5[13][45] = 4'h0;
    SS5[14][45] = 4'h0;
    SS5[15][45] = 4'h0;
    SS5[16][45] = 4'h0;
    SS5[17][45] = 4'h0;
    SS5[18][45] = 4'h0;
    SS5[19][45] = 4'h0;
    SS5[20][45] = 4'h0;
    SS5[21][45] = 4'h0;
    SS5[22][45] = 4'h0;
    SS5[23][45] = 4'h0;
    SS5[24][45] = 4'h0;
    SS5[25][45] = 4'h0;
    SS5[26][45] = 4'h0;
    SS5[27][45] = 4'h0;
    SS5[28][45] = 4'h0;
    SS5[29][45] = 4'h0;
    SS5[30][45] = 4'h0;
    SS5[31][45] = 4'h0;
    SS5[32][45] = 4'h0;
    SS5[33][45] = 4'h0;
    SS5[34][45] = 4'h0;
    SS5[35][45] = 4'h0;
    SS5[36][45] = 4'h0;
    SS5[37][45] = 4'h0;
    SS5[38][45] = 4'h0;
    SS5[39][45] = 4'h0;
    SS5[40][45] = 4'h0;
    SS5[41][45] = 4'h0;
    SS5[42][45] = 4'h0;
    SS5[43][45] = 4'h0;
    SS5[44][45] = 4'h0;
    SS5[45][45] = 4'h0;
    SS5[46][45] = 4'h0;
    SS5[47][45] = 4'h0;
    SS5[0][46] = 4'h0;
    SS5[1][46] = 4'h0;
    SS5[2][46] = 4'h0;
    SS5[3][46] = 4'h0;
    SS5[4][46] = 4'h0;
    SS5[5][46] = 4'h0;
    SS5[6][46] = 4'h0;
    SS5[7][46] = 4'h0;
    SS5[8][46] = 4'h0;
    SS5[9][46] = 4'h0;
    SS5[10][46] = 4'h0;
    SS5[11][46] = 4'h0;
    SS5[12][46] = 4'h0;
    SS5[13][46] = 4'h0;
    SS5[14][46] = 4'h0;
    SS5[15][46] = 4'h0;
    SS5[16][46] = 4'h0;
    SS5[17][46] = 4'h0;
    SS5[18][46] = 4'h0;
    SS5[19][46] = 4'h0;
    SS5[20][46] = 4'h0;
    SS5[21][46] = 4'h0;
    SS5[22][46] = 4'h0;
    SS5[23][46] = 4'h0;
    SS5[24][46] = 4'h0;
    SS5[25][46] = 4'h0;
    SS5[26][46] = 4'h0;
    SS5[27][46] = 4'h0;
    SS5[28][46] = 4'h0;
    SS5[29][46] = 4'h0;
    SS5[30][46] = 4'h0;
    SS5[31][46] = 4'h0;
    SS5[32][46] = 4'h0;
    SS5[33][46] = 4'h0;
    SS5[34][46] = 4'h0;
    SS5[35][46] = 4'h0;
    SS5[36][46] = 4'h0;
    SS5[37][46] = 4'h0;
    SS5[38][46] = 4'h0;
    SS5[39][46] = 4'h0;
    SS5[40][46] = 4'h0;
    SS5[41][46] = 4'h0;
    SS5[42][46] = 4'h0;
    SS5[43][46] = 4'h0;
    SS5[44][46] = 4'h0;
    SS5[45][46] = 4'h0;
    SS5[46][46] = 4'h0;
    SS5[47][46] = 4'h0;
    SS5[0][47] = 4'h0;
    SS5[1][47] = 4'h0;
    SS5[2][47] = 4'h0;
    SS5[3][47] = 4'h0;
    SS5[4][47] = 4'h0;
    SS5[5][47] = 4'h0;
    SS5[6][47] = 4'h0;
    SS5[7][47] = 4'h0;
    SS5[8][47] = 4'h0;
    SS5[9][47] = 4'h0;
    SS5[10][47] = 4'h0;
    SS5[11][47] = 4'h0;
    SS5[12][47] = 4'h0;
    SS5[13][47] = 4'h0;
    SS5[14][47] = 4'h0;
    SS5[15][47] = 4'h0;
    SS5[16][47] = 4'h0;
    SS5[17][47] = 4'h0;
    SS5[18][47] = 4'h0;
    SS5[19][47] = 4'h0;
    SS5[20][47] = 4'h0;
    SS5[21][47] = 4'h0;
    SS5[22][47] = 4'h0;
    SS5[23][47] = 4'h0;
    SS5[24][47] = 4'h0;
    SS5[25][47] = 4'h0;
    SS5[26][47] = 4'h0;
    SS5[27][47] = 4'h0;
    SS5[28][47] = 4'h0;
    SS5[29][47] = 4'h0;
    SS5[30][47] = 4'h0;
    SS5[31][47] = 4'h0;
    SS5[32][47] = 4'h0;
    SS5[33][47] = 4'h0;
    SS5[34][47] = 4'h0;
    SS5[35][47] = 4'h0;
    SS5[36][47] = 4'h0;
    SS5[37][47] = 4'h0;
    SS5[38][47] = 4'h0;
    SS5[39][47] = 4'h0;
    SS5[40][47] = 4'h0;
    SS5[41][47] = 4'h0;
    SS5[42][47] = 4'h0;
    SS5[43][47] = 4'h0;
    SS5[44][47] = 4'h0;
    SS5[45][47] = 4'h0;
    SS5[46][47] = 4'h0;
    SS5[47][47] = 4'h0;
 
//SS 6
    SS6[0][0] = 4'h0;
    SS6[1][0] = 4'h0;
    SS6[2][0] = 4'h0;
    SS6[3][0] = 4'h0;
    SS6[4][0] = 4'h0;
    SS6[5][0] = 4'h0;
    SS6[6][0] = 4'h0;
    SS6[7][0] = 4'h0;
    SS6[8][0] = 4'h0;
    SS6[9][0] = 4'h0;
    SS6[10][0] = 4'h0;
    SS6[11][0] = 4'h0;
    SS6[12][0] = 4'h0;
    SS6[13][0] = 4'h0;
    SS6[14][0] = 4'h0;
    SS6[15][0] = 4'h0;
    SS6[16][0] = 4'h0;
    SS6[17][0] = 4'hE;
    SS6[18][0] = 4'hC;
    SS6[19][0] = 4'hC;
    SS6[20][0] = 4'hC;
    SS6[21][0] = 4'hC;
    SS6[22][0] = 4'h0;
    SS6[23][0] = 4'h0;
    SS6[24][0] = 4'h0;
    SS6[25][0] = 4'h0;
    SS6[26][0] = 4'h0;
    SS6[27][0] = 4'h0;
    SS6[28][0] = 4'h0;
    SS6[29][0] = 4'h0;
    SS6[30][0] = 4'h0;
    SS6[31][0] = 4'h0;
    SS6[32][0] = 4'h0;
    SS6[33][0] = 4'h0;
    SS6[34][0] = 4'h0;
    SS6[35][0] = 4'h0;
    SS6[36][0] = 4'h0;
    SS6[37][0] = 4'h0;
    SS6[38][0] = 4'h0;
    SS6[39][0] = 4'h0;
    SS6[40][0] = 4'h0;
    SS6[41][0] = 4'h0;
    SS6[42][0] = 4'h0;
    SS6[43][0] = 4'h0;
    SS6[44][0] = 4'h0;
    SS6[45][0] = 4'h0;
    SS6[46][0] = 4'h0;
    SS6[47][0] = 4'h0;
    SS6[0][1] = 4'h0;
    SS6[1][1] = 4'h0;
    SS6[2][1] = 4'h0;
    SS6[3][1] = 4'h0;
    SS6[4][1] = 4'h0;
    SS6[5][1] = 4'h0;
    SS6[6][1] = 4'h0;
    SS6[7][1] = 4'h0;
    SS6[8][1] = 4'h0;
    SS6[9][1] = 4'h0;
    SS6[10][1] = 4'h0;
    SS6[11][1] = 4'h0;
    SS6[12][1] = 4'h0;
    SS6[13][1] = 4'h0;
    SS6[14][1] = 4'h0;
    SS6[15][1] = 4'h0;
    SS6[16][1] = 4'h0;
    SS6[17][1] = 4'hD;
    SS6[18][1] = 4'hC;
    SS6[19][1] = 4'hC;
    SS6[20][1] = 4'hC;
    SS6[21][1] = 4'hC;
    SS6[22][1] = 4'hC;
    SS6[23][1] = 4'h0;
    SS6[24][1] = 4'h0;
    SS6[25][1] = 4'h0;
    SS6[26][1] = 4'h0;
    SS6[27][1] = 4'h0;
    SS6[28][1] = 4'h0;
    SS6[29][1] = 4'h0;
    SS6[30][1] = 4'h0;
    SS6[31][1] = 4'h0;
    SS6[32][1] = 4'h0;
    SS6[33][1] = 4'h0;
    SS6[34][1] = 4'hD;
    SS6[35][1] = 4'h0;
    SS6[36][1] = 4'h0;
    SS6[37][1] = 4'h0;
    SS6[38][1] = 4'h0;
    SS6[39][1] = 4'h0;
    SS6[40][1] = 4'h0;
    SS6[41][1] = 4'h0;
    SS6[42][1] = 4'h0;
    SS6[43][1] = 4'h0;
    SS6[44][1] = 4'h0;
    SS6[45][1] = 4'h0;
    SS6[46][1] = 4'h0;
    SS6[47][1] = 4'h0;
    SS6[0][2] = 4'h0;
    SS6[1][2] = 4'h0;
    SS6[2][2] = 4'h0;
    SS6[3][2] = 4'h0;
    SS6[4][2] = 4'h0;
    SS6[5][2] = 4'h0;
    SS6[6][2] = 4'h0;
    SS6[7][2] = 4'h0;
    SS6[8][2] = 4'h0;
    SS6[9][2] = 4'h0;
    SS6[10][2] = 4'h0;
    SS6[11][2] = 4'h0;
    SS6[12][2] = 4'h0;
    SS6[13][2] = 4'h0;
    SS6[14][2] = 4'h0;
    SS6[15][2] = 4'h0;
    SS6[16][2] = 4'hD;
    SS6[17][2] = 4'hD;
    SS6[18][2] = 4'hD;
    SS6[19][2] = 4'hC;
    SS6[20][2] = 4'hC;
    SS6[21][2] = 4'hC;
    SS6[22][2] = 4'hC;
    SS6[23][2] = 4'hC;
    SS6[24][2] = 4'h0;
    SS6[25][2] = 4'h0;
    SS6[26][2] = 4'h0;
    SS6[27][2] = 4'h0;
    SS6[28][2] = 4'h0;
    SS6[29][2] = 4'h0;
    SS6[30][2] = 4'h0;
    SS6[31][2] = 4'h0;
    SS6[32][2] = 4'h0;
    SS6[33][2] = 4'hD;
    SS6[34][2] = 4'hD;
    SS6[35][2] = 4'hD;
    SS6[36][2] = 4'h0;
    SS6[37][2] = 4'h0;
    SS6[38][2] = 4'h0;
    SS6[39][2] = 4'h0;
    SS6[40][2] = 4'h0;
    SS6[41][2] = 4'h0;
    SS6[42][2] = 4'h0;
    SS6[43][2] = 4'h0;
    SS6[44][2] = 4'h0;
    SS6[45][2] = 4'h0;
    SS6[46][2] = 4'h0;
    SS6[47][2] = 4'h0;
    SS6[0][3] = 4'h0;
    SS6[1][3] = 4'h0;
    SS6[2][3] = 4'h0;
    SS6[3][3] = 4'h0;
    SS6[4][3] = 4'h0;
    SS6[5][3] = 4'h0;
    SS6[6][3] = 4'h0;
    SS6[7][3] = 4'h0;
    SS6[8][3] = 4'h0;
    SS6[9][3] = 4'h0;
    SS6[10][3] = 4'h0;
    SS6[11][3] = 4'h0;
    SS6[12][3] = 4'h0;
    SS6[13][3] = 4'h0;
    SS6[14][3] = 4'h0;
    SS6[15][3] = 4'h0;
    SS6[16][3] = 4'hD;
    SS6[17][3] = 4'hD;
    SS6[18][3] = 4'hD;
    SS6[19][3] = 4'hC;
    SS6[20][3] = 4'hC;
    SS6[21][3] = 4'hC;
    SS6[22][3] = 4'hC;
    SS6[23][3] = 4'h0;
    SS6[24][3] = 4'h0;
    SS6[25][3] = 4'h0;
    SS6[26][3] = 4'h0;
    SS6[27][3] = 4'h0;
    SS6[28][3] = 4'h0;
    SS6[29][3] = 4'h0;
    SS6[30][3] = 4'h0;
    SS6[31][3] = 4'h0;
    SS6[32][3] = 4'hD;
    SS6[33][3] = 4'hD;
    SS6[34][3] = 4'hD;
    SS6[35][3] = 4'hD;
    SS6[36][3] = 4'h0;
    SS6[37][3] = 4'h0;
    SS6[38][3] = 4'h0;
    SS6[39][3] = 4'h0;
    SS6[40][3] = 4'h0;
    SS6[41][3] = 4'h0;
    SS6[42][3] = 4'h0;
    SS6[43][3] = 4'h0;
    SS6[44][3] = 4'h0;
    SS6[45][3] = 4'h0;
    SS6[46][3] = 4'h0;
    SS6[47][3] = 4'h0;
    SS6[0][4] = 4'h0;
    SS6[1][4] = 4'h0;
    SS6[2][4] = 4'h0;
    SS6[3][4] = 4'h0;
    SS6[4][4] = 4'h0;
    SS6[5][4] = 4'h0;
    SS6[6][4] = 4'h0;
    SS6[7][4] = 4'h0;
    SS6[8][4] = 4'h0;
    SS6[9][4] = 4'h0;
    SS6[10][4] = 4'h0;
    SS6[11][4] = 4'h0;
    SS6[12][4] = 4'h0;
    SS6[13][4] = 4'h0;
    SS6[14][4] = 4'h0;
    SS6[15][4] = 4'h0;
    SS6[16][4] = 4'h0;
    SS6[17][4] = 4'hD;
    SS6[18][4] = 4'hC;
    SS6[19][4] = 4'hC;
    SS6[20][4] = 4'hC;
    SS6[21][4] = 4'hC;
    SS6[22][4] = 4'h0;
    SS6[23][4] = 4'h0;
    SS6[24][4] = 4'h0;
    SS6[25][4] = 4'h0;
    SS6[26][4] = 4'h0;
    SS6[27][4] = 4'h0;
    SS6[28][4] = 4'h0;
    SS6[29][4] = 4'h0;
    SS6[30][4] = 4'h0;
    SS6[31][4] = 4'hD;
    SS6[32][4] = 4'hD;
    SS6[33][4] = 4'hD;
    SS6[34][4] = 4'hD;
    SS6[35][4] = 4'h0;
    SS6[36][4] = 4'h0;
    SS6[37][4] = 4'h0;
    SS6[38][4] = 4'h0;
    SS6[39][4] = 4'h0;
    SS6[40][4] = 4'h0;
    SS6[41][4] = 4'h0;
    SS6[42][4] = 4'h0;
    SS6[43][4] = 4'h0;
    SS6[44][4] = 4'h0;
    SS6[45][4] = 4'h0;
    SS6[46][4] = 4'h0;
    SS6[47][4] = 4'h0;
    SS6[0][5] = 4'h0;
    SS6[1][5] = 4'h0;
    SS6[2][5] = 4'h0;
    SS6[3][5] = 4'h0;
    SS6[4][5] = 4'h0;
    SS6[5][5] = 4'h0;
    SS6[6][5] = 4'h0;
    SS6[7][5] = 4'h0;
    SS6[8][5] = 4'h0;
    SS6[9][5] = 4'h0;
    SS6[10][5] = 4'h0;
    SS6[11][5] = 4'h0;
    SS6[12][5] = 4'h0;
    SS6[13][5] = 4'h0;
    SS6[14][5] = 4'h0;
    SS6[15][5] = 4'h0;
    SS6[16][5] = 4'h0;
    SS6[17][5] = 4'hE;
    SS6[18][5] = 4'hC;
    SS6[19][5] = 4'hC;
    SS6[20][5] = 4'hC;
    SS6[21][5] = 4'hC;
    SS6[22][5] = 4'h0;
    SS6[23][5] = 4'h0;
    SS6[24][5] = 4'h0;
    SS6[25][5] = 4'h0;
    SS6[26][5] = 4'h0;
    SS6[27][5] = 4'h0;
    SS6[28][5] = 4'h0;
    SS6[29][5] = 4'h0;
    SS6[30][5] = 4'hE;
    SS6[31][5] = 4'hD;
    SS6[32][5] = 4'hD;
    SS6[33][5] = 4'hD;
    SS6[34][5] = 4'hD;
    SS6[35][5] = 4'h0;
    SS6[36][5] = 4'h0;
    SS6[37][5] = 4'h0;
    SS6[38][5] = 4'h0;
    SS6[39][5] = 4'h0;
    SS6[40][5] = 4'h0;
    SS6[41][5] = 4'h0;
    SS6[42][5] = 4'h0;
    SS6[43][5] = 4'h0;
    SS6[44][5] = 4'h0;
    SS6[45][5] = 4'h0;
    SS6[46][5] = 4'h0;
    SS6[47][5] = 4'h0;
    SS6[0][6] = 4'h0;
    SS6[1][6] = 4'h0;
    SS6[2][6] = 4'h0;
    SS6[3][6] = 4'h0;
    SS6[4][6] = 4'h0;
    SS6[5][6] = 4'h0;
    SS6[6][6] = 4'h0;
    SS6[7][6] = 4'h0;
    SS6[8][6] = 4'h0;
    SS6[9][6] = 4'h0;
    SS6[10][6] = 4'h0;
    SS6[11][6] = 4'h0;
    SS6[12][6] = 4'h0;
    SS6[13][6] = 4'h0;
    SS6[14][6] = 4'h0;
    SS6[15][6] = 4'h0;
    SS6[16][6] = 4'hE;
    SS6[17][6] = 4'hE;
    SS6[18][6] = 4'hE;
    SS6[19][6] = 4'hC;
    SS6[20][6] = 4'hC;
    SS6[21][6] = 4'hC;
    SS6[22][6] = 4'hC;
    SS6[23][6] = 4'h0;
    SS6[24][6] = 4'h0;
    SS6[25][6] = 4'h0;
    SS6[26][6] = 4'h0;
    SS6[27][6] = 4'h0;
    SS6[28][6] = 4'h0;
    SS6[29][6] = 4'hE;
    SS6[30][6] = 4'hE;
    SS6[31][6] = 4'hE;
    SS6[32][6] = 4'hD;
    SS6[33][6] = 4'hD;
    SS6[34][6] = 4'hD;
    SS6[35][6] = 4'hD;
    SS6[36][6] = 4'h0;
    SS6[37][6] = 4'h0;
    SS6[38][6] = 4'h0;
    SS6[39][6] = 4'h0;
    SS6[40][6] = 4'h0;
    SS6[41][6] = 4'h0;
    SS6[42][6] = 4'h0;
    SS6[43][6] = 4'h0;
    SS6[44][6] = 4'h0;
    SS6[45][6] = 4'h0;
    SS6[46][6] = 4'h0;
    SS6[47][6] = 4'h0;
    SS6[0][7] = 4'h0;
    SS6[1][7] = 4'h0;
    SS6[2][7] = 4'h0;
    SS6[3][7] = 4'h0;
    SS6[4][7] = 4'h0;
    SS6[5][7] = 4'h0;
    SS6[6][7] = 4'h0;
    SS6[7][7] = 4'h0;
    SS6[8][7] = 4'h0;
    SS6[9][7] = 4'h0;
    SS6[10][7] = 4'h0;
    SS6[11][7] = 4'h0;
    SS6[12][7] = 4'h0;
    SS6[13][7] = 4'h0;
    SS6[14][7] = 4'h0;
    SS6[15][7] = 4'h0;
    SS6[16][7] = 4'hE;
    SS6[17][7] = 4'hE;
    SS6[18][7] = 4'hE;
    SS6[19][7] = 4'hD;
    SS6[20][7] = 4'hC;
    SS6[21][7] = 4'hC;
    SS6[22][7] = 4'hC;
    SS6[23][7] = 4'hC;
    SS6[24][7] = 4'hD;
    SS6[25][7] = 4'h0;
    SS6[26][7] = 4'h0;
    SS6[27][7] = 4'h0;
    SS6[28][7] = 4'hE;
    SS6[29][7] = 4'hE;
    SS6[30][7] = 4'hE;
    SS6[31][7] = 4'hE;
    SS6[32][7] = 4'hD;
    SS6[33][7] = 4'hD;
    SS6[34][7] = 4'hD;
    SS6[35][7] = 4'hD;
    SS6[36][7] = 4'h0;
    SS6[37][7] = 4'h0;
    SS6[38][7] = 4'h0;
    SS6[39][7] = 4'h0;
    SS6[40][7] = 4'h0;
    SS6[41][7] = 4'h0;
    SS6[42][7] = 4'h0;
    SS6[43][7] = 4'h0;
    SS6[44][7] = 4'h0;
    SS6[45][7] = 4'h0;
    SS6[46][7] = 4'h0;
    SS6[47][7] = 4'h0;
    SS6[0][8] = 4'h0;
    SS6[1][8] = 4'h0;
    SS6[2][8] = 4'h0;
    SS6[3][8] = 4'h0;
    SS6[4][8] = 4'h0;
    SS6[5][8] = 4'h0;
    SS6[6][8] = 4'h0;
    SS6[7][8] = 4'h0;
    SS6[8][8] = 4'h0;
    SS6[9][8] = 4'h0;
    SS6[10][8] = 4'h0;
    SS6[11][8] = 4'h0;
    SS6[12][8] = 4'h0;
    SS6[13][8] = 4'h0;
    SS6[14][8] = 4'h0;
    SS6[15][8] = 4'h0;
    SS6[16][8] = 4'h0;
    SS6[17][8] = 4'hE;
    SS6[18][8] = 4'hD;
    SS6[19][8] = 4'hD;
    SS6[20][8] = 4'hD;
    SS6[21][8] = 4'hC;
    SS6[22][8] = 4'hC;
    SS6[23][8] = 4'hC;
    SS6[24][8] = 4'hC;
    SS6[25][8] = 4'hD;
    SS6[26][8] = 4'h0;
    SS6[27][8] = 4'hE;
    SS6[28][8] = 4'hE;
    SS6[29][8] = 4'hE;
    SS6[30][8] = 4'hE;
    SS6[31][8] = 4'hD;
    SS6[32][8] = 4'hD;
    SS6[33][8] = 4'hD;
    SS6[34][8] = 4'hD;
    SS6[35][8] = 4'h0;
    SS6[36][8] = 4'h0;
    SS6[37][8] = 4'h0;
    SS6[38][8] = 4'h0;
    SS6[39][8] = 4'h0;
    SS6[40][8] = 4'h0;
    SS6[41][8] = 4'h0;
    SS6[42][8] = 4'h0;
    SS6[43][8] = 4'h0;
    SS6[44][8] = 4'h0;
    SS6[45][8] = 4'h0;
    SS6[46][8] = 4'h0;
    SS6[47][8] = 4'h0;
    SS6[0][9] = 4'h0;
    SS6[1][9] = 4'h0;
    SS6[2][9] = 4'h0;
    SS6[3][9] = 4'h0;
    SS6[4][9] = 4'h0;
    SS6[5][9] = 4'h0;
    SS6[6][9] = 4'h0;
    SS6[7][9] = 4'h0;
    SS6[8][9] = 4'h0;
    SS6[9][9] = 4'h0;
    SS6[10][9] = 4'h0;
    SS6[11][9] = 4'h0;
    SS6[12][9] = 4'h0;
    SS6[13][9] = 4'h0;
    SS6[14][9] = 4'h0;
    SS6[15][9] = 4'h0;
    SS6[16][9] = 4'h0;
    SS6[17][9] = 4'hE;
    SS6[18][9] = 4'hD;
    SS6[19][9] = 4'hD;
    SS6[20][9] = 4'hD;
    SS6[21][9] = 4'hD;
    SS6[22][9] = 4'hC;
    SS6[23][9] = 4'hC;
    SS6[24][9] = 4'hC;
    SS6[25][9] = 4'hC;
    SS6[26][9] = 4'hE;
    SS6[27][9] = 4'hE;
    SS6[28][9] = 4'hE;
    SS6[29][9] = 4'hE;
    SS6[30][9] = 4'hE;
    SS6[31][9] = 4'hD;
    SS6[32][9] = 4'hD;
    SS6[33][9] = 4'hD;
    SS6[34][9] = 4'h3;
    SS6[35][9] = 4'h0;
    SS6[36][9] = 4'h0;
    SS6[37][9] = 4'h0;
    SS6[38][9] = 4'h0;
    SS6[39][9] = 4'h0;
    SS6[40][9] = 4'h0;
    SS6[41][9] = 4'h0;
    SS6[42][9] = 4'h0;
    SS6[43][9] = 4'h0;
    SS6[44][9] = 4'h0;
    SS6[45][9] = 4'h0;
    SS6[46][9] = 4'h0;
    SS6[47][9] = 4'h0;
    SS6[0][10] = 4'h0;
    SS6[1][10] = 4'h0;
    SS6[2][10] = 4'h0;
    SS6[3][10] = 4'h0;
    SS6[4][10] = 4'h0;
    SS6[5][10] = 4'h0;
    SS6[6][10] = 4'h0;
    SS6[7][10] = 4'h0;
    SS6[8][10] = 4'h0;
    SS6[9][10] = 4'h0;
    SS6[10][10] = 4'h0;
    SS6[11][10] = 4'h0;
    SS6[12][10] = 4'h0;
    SS6[13][10] = 4'h0;
    SS6[14][10] = 4'h0;
    SS6[15][10] = 4'h0;
    SS6[16][10] = 4'hE;
    SS6[17][10] = 4'hE;
    SS6[18][10] = 4'hE;
    SS6[19][10] = 4'hD;
    SS6[20][10] = 4'hD;
    SS6[21][10] = 4'hC;
    SS6[22][10] = 4'hC;
    SS6[23][10] = 4'hC;
    SS6[24][10] = 4'hC;
    SS6[25][10] = 4'hC;
    SS6[26][10] = 4'hC;
    SS6[27][10] = 4'hE;
    SS6[28][10] = 4'hE;
    SS6[29][10] = 4'hE;
    SS6[30][10] = 4'hE;
    SS6[31][10] = 4'hE;
    SS6[32][10] = 4'hD;
    SS6[33][10] = 4'h3;
    SS6[34][10] = 4'h3;
    SS6[35][10] = 4'h3;
    SS6[36][10] = 4'h0;
    SS6[37][10] = 4'h0;
    SS6[38][10] = 4'h0;
    SS6[39][10] = 4'h0;
    SS6[40][10] = 4'h0;
    SS6[41][10] = 4'h0;
    SS6[42][10] = 4'h0;
    SS6[43][10] = 4'h0;
    SS6[44][10] = 4'h0;
    SS6[45][10] = 4'h0;
    SS6[46][10] = 4'h0;
    SS6[47][10] = 4'h0;
    SS6[0][11] = 4'h0;
    SS6[1][11] = 4'h0;
    SS6[2][11] = 4'h0;
    SS6[3][11] = 4'h0;
    SS6[4][11] = 4'h0;
    SS6[5][11] = 4'h0;
    SS6[6][11] = 4'h0;
    SS6[7][11] = 4'h0;
    SS6[8][11] = 4'h0;
    SS6[9][11] = 4'h0;
    SS6[10][11] = 4'h0;
    SS6[11][11] = 4'h0;
    SS6[12][11] = 4'h0;
    SS6[13][11] = 4'h0;
    SS6[14][11] = 4'h0;
    SS6[15][11] = 4'h0;
    SS6[16][11] = 4'hE;
    SS6[17][11] = 4'hE;
    SS6[18][11] = 4'hE;
    SS6[19][11] = 4'hD;
    SS6[20][11] = 4'hC;
    SS6[21][11] = 4'hC;
    SS6[22][11] = 4'hC;
    SS6[23][11] = 4'hC;
    SS6[24][11] = 4'hC;
    SS6[25][11] = 4'hC;
    SS6[26][11] = 4'hC;
    SS6[27][11] = 4'hC;
    SS6[28][11] = 4'hE;
    SS6[29][11] = 4'hE;
    SS6[30][11] = 4'hE;
    SS6[31][11] = 4'hE;
    SS6[32][11] = 4'hD;
    SS6[33][11] = 4'h3;
    SS6[34][11] = 4'h3;
    SS6[35][11] = 4'h3;
    SS6[36][11] = 4'h2;
    SS6[37][11] = 4'h0;
    SS6[38][11] = 4'h0;
    SS6[39][11] = 4'h0;
    SS6[40][11] = 4'h0;
    SS6[41][11] = 4'h0;
    SS6[42][11] = 4'h0;
    SS6[43][11] = 4'h0;
    SS6[44][11] = 4'h0;
    SS6[45][11] = 4'h0;
    SS6[46][11] = 4'h0;
    SS6[47][11] = 4'h0;
    SS6[0][12] = 4'h0;
    SS6[1][12] = 4'h0;
    SS6[2][12] = 4'h0;
    SS6[3][12] = 4'h0;
    SS6[4][12] = 4'h0;
    SS6[5][12] = 4'h0;
    SS6[6][12] = 4'h0;
    SS6[7][12] = 4'h0;
    SS6[8][12] = 4'h0;
    SS6[9][12] = 4'h0;
    SS6[10][12] = 4'h0;
    SS6[11][12] = 4'h0;
    SS6[12][12] = 4'h0;
    SS6[13][12] = 4'h0;
    SS6[14][12] = 4'h0;
    SS6[15][12] = 4'h0;
    SS6[16][12] = 4'h0;
    SS6[17][12] = 4'hE;
    SS6[18][12] = 4'hD;
    SS6[19][12] = 4'hD;
    SS6[20][12] = 4'hD;
    SS6[21][12] = 4'hC;
    SS6[22][12] = 4'hC;
    SS6[23][12] = 4'hC;
    SS6[24][12] = 4'hC;
    SS6[25][12] = 4'hC;
    SS6[26][12] = 4'hC;
    SS6[27][12] = 4'hE;
    SS6[28][12] = 4'hE;
    SS6[29][12] = 4'hE;
    SS6[30][12] = 4'hE;
    SS6[31][12] = 4'hD;
    SS6[32][12] = 4'hD;
    SS6[33][12] = 4'hD;
    SS6[34][12] = 4'h3;
    SS6[35][12] = 4'h2;
    SS6[36][12] = 4'h0;
    SS6[37][12] = 4'h0;
    SS6[38][12] = 4'h0;
    SS6[39][12] = 4'h0;
    SS6[40][12] = 4'h0;
    SS6[41][12] = 4'h0;
    SS6[42][12] = 4'h0;
    SS6[43][12] = 4'h0;
    SS6[44][12] = 4'h0;
    SS6[45][12] = 4'h0;
    SS6[46][12] = 4'h0;
    SS6[47][12] = 4'h0;
    SS6[0][13] = 4'h0;
    SS6[1][13] = 4'h0;
    SS6[2][13] = 4'h0;
    SS6[3][13] = 4'h0;
    SS6[4][13] = 4'h0;
    SS6[5][13] = 4'h0;
    SS6[6][13] = 4'h0;
    SS6[7][13] = 4'h0;
    SS6[8][13] = 4'h0;
    SS6[9][13] = 4'h0;
    SS6[10][13] = 4'h0;
    SS6[11][13] = 4'h0;
    SS6[12][13] = 4'h0;
    SS6[13][13] = 4'h0;
    SS6[14][13] = 4'h0;
    SS6[15][13] = 4'h0;
    SS6[16][13] = 4'h0;
    SS6[17][13] = 4'h0;
    SS6[18][13] = 4'hD;
    SS6[19][13] = 4'hD;
    SS6[20][13] = 4'hD;
    SS6[21][13] = 4'hD;
    SS6[22][13] = 4'hC;
    SS6[23][13] = 4'hC;
    SS6[24][13] = 4'hC;
    SS6[25][13] = 4'hC;
    SS6[26][13] = 4'hE;
    SS6[27][13] = 4'hE;
    SS6[28][13] = 4'hE;
    SS6[29][13] = 4'hE;
    SS6[30][13] = 4'hD;
    SS6[31][13] = 4'hD;
    SS6[32][13] = 4'hD;
    SS6[33][13] = 4'hD;
    SS6[34][13] = 4'hE;
    SS6[35][13] = 4'h0;
    SS6[36][13] = 4'h0;
    SS6[37][13] = 4'h0;
    SS6[38][13] = 4'h0;
    SS6[39][13] = 4'h0;
    SS6[40][13] = 4'h0;
    SS6[41][13] = 4'h0;
    SS6[42][13] = 4'h0;
    SS6[43][13] = 4'h0;
    SS6[44][13] = 4'h0;
    SS6[45][13] = 4'h0;
    SS6[46][13] = 4'h0;
    SS6[47][13] = 4'h0;
    SS6[0][14] = 4'h0;
    SS6[1][14] = 4'h0;
    SS6[2][14] = 4'h0;
    SS6[3][14] = 4'h0;
    SS6[4][14] = 4'h0;
    SS6[5][14] = 4'h0;
    SS6[6][14] = 4'h0;
    SS6[7][14] = 4'h0;
    SS6[8][14] = 4'h0;
    SS6[9][14] = 4'h0;
    SS6[10][14] = 4'h0;
    SS6[11][14] = 4'h0;
    SS6[12][14] = 4'h0;
    SS6[13][14] = 4'h0;
    SS6[14][14] = 4'h0;
    SS6[15][14] = 4'h0;
    SS6[16][14] = 4'h0;
    SS6[17][14] = 4'hE;
    SS6[18][14] = 4'hE;
    SS6[19][14] = 4'hD;
    SS6[20][14] = 4'hD;
    SS6[21][14] = 4'hC;
    SS6[22][14] = 4'hC;
    SS6[23][14] = 4'hC;
    SS6[24][14] = 4'hC;
    SS6[25][14] = 4'hC;
    SS6[26][14] = 4'hC;
    SS6[27][14] = 4'hE;
    SS6[28][14] = 4'hE;
    SS6[29][14] = 4'hD;
    SS6[30][14] = 4'hD;
    SS6[31][14] = 4'hD;
    SS6[32][14] = 4'hD;
    SS6[33][14] = 4'hE;
    SS6[34][14] = 4'h0;
    SS6[35][14] = 4'h0;
    SS6[36][14] = 4'h0;
    SS6[37][14] = 4'h0;
    SS6[38][14] = 4'h0;
    SS6[39][14] = 4'h0;
    SS6[40][14] = 4'h0;
    SS6[41][14] = 4'h0;
    SS6[42][14] = 4'h0;
    SS6[43][14] = 4'h0;
    SS6[44][14] = 4'h0;
    SS6[45][14] = 4'h0;
    SS6[46][14] = 4'h0;
    SS6[47][14] = 4'h0;
    SS6[0][15] = 4'h0;
    SS6[1][15] = 4'h0;
    SS6[2][15] = 4'h0;
    SS6[3][15] = 4'h0;
    SS6[4][15] = 4'h0;
    SS6[5][15] = 4'h0;
    SS6[6][15] = 4'h0;
    SS6[7][15] = 4'h0;
    SS6[8][15] = 4'h0;
    SS6[9][15] = 4'h0;
    SS6[10][15] = 4'h0;
    SS6[11][15] = 4'h0;
    SS6[12][15] = 4'h0;
    SS6[13][15] = 4'h0;
    SS6[14][15] = 4'h0;
    SS6[15][15] = 4'hF;
    SS6[16][15] = 4'hE;
    SS6[17][15] = 4'hE;
    SS6[18][15] = 4'hE;
    SS6[19][15] = 4'hE;
    SS6[20][15] = 4'hC;
    SS6[21][15] = 4'hC;
    SS6[22][15] = 4'hC;
    SS6[23][15] = 4'hC;
    SS6[24][15] = 4'hC;
    SS6[25][15] = 4'hC;
    SS6[26][15] = 4'hC;
    SS6[27][15] = 4'hC;
    SS6[28][15] = 4'hD;
    SS6[29][15] = 4'hD;
    SS6[30][15] = 4'hD;
    SS6[31][15] = 4'hD;
    SS6[32][15] = 4'hD;
    SS6[33][15] = 4'h0;
    SS6[34][15] = 4'h0;
    SS6[35][15] = 4'h0;
    SS6[36][15] = 4'h0;
    SS6[37][15] = 4'h0;
    SS6[38][15] = 4'h0;
    SS6[39][15] = 4'h0;
    SS6[40][15] = 4'h0;
    SS6[41][15] = 4'h0;
    SS6[42][15] = 4'h0;
    SS6[43][15] = 4'h0;
    SS6[44][15] = 4'h0;
    SS6[45][15] = 4'h0;
    SS6[46][15] = 4'h0;
    SS6[47][15] = 4'h0;
    SS6[0][16] = 4'h0;
    SS6[1][16] = 4'h0;
    SS6[2][16] = 4'hD;
    SS6[3][16] = 4'hD;
    SS6[4][16] = 4'h0;
    SS6[5][16] = 4'h0;
    SS6[6][16] = 4'hE;
    SS6[7][16] = 4'hE;
    SS6[8][16] = 4'h0;
    SS6[9][16] = 4'h0;
    SS6[10][16] = 4'hE;
    SS6[11][16] = 4'hE;
    SS6[12][16] = 4'h0;
    SS6[13][16] = 4'h0;
    SS6[14][16] = 4'h0;
    SS6[15][16] = 4'hE;
    SS6[16][16] = 4'hE;
    SS6[17][16] = 4'hE;
    SS6[18][16] = 4'hE;
    SS6[19][16] = 4'hE;
    SS6[20][16] = 4'hE;
    SS6[21][16] = 4'hC;
    SS6[22][16] = 4'hC;
    SS6[23][16] = 4'hC;
    SS6[24][16] = 4'hC;
    SS6[25][16] = 4'hC;
    SS6[26][16] = 4'hC;
    SS6[27][16] = 4'hE;
    SS6[28][16] = 4'hE;
    SS6[29][16] = 4'hD;
    SS6[30][16] = 4'hD;
    SS6[31][16] = 4'hD;
    SS6[32][16] = 4'hD;
    SS6[33][16] = 4'h0;
    SS6[34][16] = 4'h0;
    SS6[35][16] = 4'h0;
    SS6[36][16] = 4'h0;
    SS6[37][16] = 4'h0;
    SS6[38][16] = 4'h0;
    SS6[39][16] = 4'h0;
    SS6[40][16] = 4'h0;
    SS6[41][16] = 4'h0;
    SS6[42][16] = 4'h0;
    SS6[43][16] = 4'h0;
    SS6[44][16] = 4'h0;
    SS6[45][16] = 4'h0;
    SS6[46][16] = 4'h0;
    SS6[47][16] = 4'h0;
    SS6[0][17] = 4'hE;
    SS6[1][17] = 4'hD;
    SS6[2][17] = 4'hD;
    SS6[3][17] = 4'hD;
    SS6[4][17] = 4'hD;
    SS6[5][17] = 4'hE;
    SS6[6][17] = 4'hE;
    SS6[7][17] = 4'hE;
    SS6[8][17] = 4'hE;
    SS6[9][17] = 4'hE;
    SS6[10][17] = 4'hE;
    SS6[11][17] = 4'hE;
    SS6[12][17] = 4'hE;
    SS6[13][17] = 4'h0;
    SS6[14][17] = 4'hE;
    SS6[15][17] = 4'hE;
    SS6[16][17] = 4'hE;
    SS6[17][17] = 4'hE;
    SS6[18][17] = 4'hE;
    SS6[19][17] = 4'hE;
    SS6[20][17] = 4'hE;
    SS6[21][17] = 4'hE;
    SS6[22][17] = 4'hC;
    SS6[23][17] = 4'hC;
    SS6[24][17] = 4'hC;
    SS6[25][17] = 4'hC;
    SS6[26][17] = 4'hE;
    SS6[27][17] = 4'hE;
    SS6[28][17] = 4'hE;
    SS6[29][17] = 4'hE;
    SS6[30][17] = 4'hD;
    SS6[31][17] = 4'hD;
    SS6[32][17] = 4'hD;
    SS6[33][17] = 4'hD;
    SS6[34][17] = 4'h0;
    SS6[35][17] = 4'h0;
    SS6[36][17] = 4'h0;
    SS6[37][17] = 4'h0;
    SS6[38][17] = 4'h0;
    SS6[39][17] = 4'h0;
    SS6[40][17] = 4'h0;
    SS6[41][17] = 4'h0;
    SS6[42][17] = 4'h0;
    SS6[43][17] = 4'h0;
    SS6[44][17] = 4'h0;
    SS6[45][17] = 4'h0;
    SS6[46][17] = 4'h0;
    SS6[47][17] = 4'h0;
    SS6[0][18] = 4'hC;
    SS6[1][18] = 4'hC;
    SS6[2][18] = 4'hD;
    SS6[3][18] = 4'hD;
    SS6[4][18] = 4'hC;
    SS6[5][18] = 4'hC;
    SS6[6][18] = 4'hE;
    SS6[7][18] = 4'hE;
    SS6[8][18] = 4'hD;
    SS6[9][18] = 4'hD;
    SS6[10][18] = 4'hE;
    SS6[11][18] = 4'hE;
    SS6[12][18] = 4'hD;
    SS6[13][18] = 4'hD;
    SS6[14][18] = 4'hE;
    SS6[15][18] = 4'hE;
    SS6[16][18] = 4'hE;
    SS6[17][18] = 4'hE;
    SS6[18][18] = 4'hE;
    SS6[19][18] = 4'hE;
    SS6[20][18] = 4'hE;
    SS6[21][18] = 4'hD;
    SS6[22][18] = 4'hD;
    SS6[23][18] = 4'hC;
    SS6[24][18] = 4'hC;
    SS6[25][18] = 4'hC;
    SS6[26][18] = 4'hC;
    SS6[27][18] = 4'hE;
    SS6[28][18] = 4'hE;
    SS6[29][18] = 4'hD;
    SS6[30][18] = 4'hD;
    SS6[31][18] = 4'hD;
    SS6[32][18] = 4'hD;
    SS6[33][18] = 4'hD;
    SS6[34][18] = 4'h3;
    SS6[35][18] = 4'h2;
    SS6[36][18] = 4'h0;
    SS6[37][18] = 4'h0;
    SS6[38][18] = 4'h0;
    SS6[39][18] = 4'h0;
    SS6[40][18] = 4'h0;
    SS6[41][18] = 4'h0;
    SS6[42][18] = 4'h0;
    SS6[43][18] = 4'h0;
    SS6[44][18] = 4'h0;
    SS6[45][18] = 4'h0;
    SS6[46][18] = 4'h0;
    SS6[47][18] = 4'h0;
    SS6[0][19] = 4'hC;
    SS6[1][19] = 4'hC;
    SS6[2][19] = 4'hC;
    SS6[3][19] = 4'hC;
    SS6[4][19] = 4'hC;
    SS6[5][19] = 4'hC;
    SS6[6][19] = 4'hC;
    SS6[7][19] = 4'hD;
    SS6[8][19] = 4'hD;
    SS6[9][19] = 4'hD;
    SS6[10][19] = 4'hD;
    SS6[11][19] = 4'hD;
    SS6[12][19] = 4'hD;
    SS6[13][19] = 4'hD;
    SS6[14][19] = 4'hD;
    SS6[15][19] = 4'hE;
    SS6[16][19] = 4'hE;
    SS6[17][19] = 4'hE;
    SS6[18][19] = 4'hE;
    SS6[19][19] = 4'hE;
    SS6[20][19] = 4'hD;
    SS6[21][19] = 4'hD;
    SS6[22][19] = 4'hD;
    SS6[23][19] = 4'hD;
    SS6[24][19] = 4'hC;
    SS6[25][19] = 4'hC;
    SS6[26][19] = 4'hC;
    SS6[27][19] = 4'hC;
    SS6[28][19] = 4'hD;
    SS6[29][19] = 4'hD;
    SS6[30][19] = 4'hD;
    SS6[31][19] = 4'hD;
    SS6[32][19] = 4'hD;
    SS6[33][19] = 4'h3;
    SS6[34][19] = 4'h3;
    SS6[35][19] = 4'h3;
    SS6[36][19] = 4'h2;
    SS6[37][19] = 4'h0;
    SS6[38][19] = 4'h0;
    SS6[39][19] = 4'h0;
    SS6[40][19] = 4'h0;
    SS6[41][19] = 4'h0;
    SS6[42][19] = 4'h0;
    SS6[43][19] = 4'h0;
    SS6[44][19] = 4'h0;
    SS6[45][19] = 4'h0;
    SS6[46][19] = 4'h0;
    SS6[47][19] = 4'h0;
    SS6[0][20] = 4'hC;
    SS6[1][20] = 4'hC;
    SS6[2][20] = 4'hC;
    SS6[3][20] = 4'hC;
    SS6[4][20] = 4'hC;
    SS6[5][20] = 4'hC;
    SS6[6][20] = 4'hC;
    SS6[7][20] = 4'hC;
    SS6[8][20] = 4'hD;
    SS6[9][20] = 4'hD;
    SS6[10][20] = 4'hD;
    SS6[11][20] = 4'hC;
    SS6[12][20] = 4'hD;
    SS6[13][20] = 4'hD;
    SS6[14][20] = 4'hD;
    SS6[15][20] = 4'hC;
    SS6[16][20] = 4'hE;
    SS6[17][20] = 4'hE;
    SS6[18][20] = 4'hE;
    SS6[19][20] = 4'hD;
    SS6[20][20] = 4'hD;
    SS6[21][20] = 4'hD;
    SS6[22][20] = 4'hD;
    SS6[23][20] = 4'hC;
    SS6[24][20] = 4'hC;
    SS6[25][20] = 4'hC;
    SS6[26][20] = 4'hC;
    SS6[27][20] = 4'hC;
    SS6[28][20] = 4'hC;
    SS6[29][20] = 4'hD;
    SS6[30][20] = 4'hD;
    SS6[31][20] = 4'hD;
    SS6[32][20] = 4'hD;
    SS6[33][20] = 4'h3;
    SS6[34][20] = 4'h3;
    SS6[35][20] = 4'h3;
    SS6[36][20] = 4'h0;
    SS6[37][20] = 4'h0;
    SS6[38][20] = 4'h0;
    SS6[39][20] = 4'h0;
    SS6[40][20] = 4'h0;
    SS6[41][20] = 4'h0;
    SS6[42][20] = 4'h0;
    SS6[43][20] = 4'h0;
    SS6[44][20] = 4'h0;
    SS6[45][20] = 4'h0;
    SS6[46][20] = 4'h0;
    SS6[47][20] = 4'h0;
    SS6[0][21] = 4'hC;
    SS6[1][21] = 4'hC;
    SS6[2][21] = 4'hC;
    SS6[3][21] = 4'hC;
    SS6[4][21] = 4'hC;
    SS6[5][21] = 4'hC;
    SS6[6][21] = 4'hC;
    SS6[7][21] = 4'hC;
    SS6[8][21] = 4'hC;
    SS6[9][21] = 4'hD;
    SS6[10][21] = 4'hC;
    SS6[11][21] = 4'hC;
    SS6[12][21] = 4'hC;
    SS6[13][21] = 4'hD;
    SS6[14][21] = 4'hC;
    SS6[15][21] = 4'hC;
    SS6[16][21] = 4'hC;
    SS6[17][21] = 4'hE;
    SS6[18][21] = 4'hD;
    SS6[19][21] = 4'hD;
    SS6[20][21] = 4'hD;
    SS6[21][21] = 4'hD;
    SS6[22][21] = 4'hC;
    SS6[23][21] = 4'hC;
    SS6[24][21] = 4'hC;
    SS6[25][21] = 4'hC;
    SS6[26][21] = 4'hC;
    SS6[27][21] = 4'hC;
    SS6[28][21] = 4'hC;
    SS6[29][21] = 4'hC;
    SS6[30][21] = 4'hD;
    SS6[31][21] = 4'hD;
    SS6[32][21] = 4'hD;
    SS6[33][21] = 4'hD;
    SS6[34][21] = 4'h3;
    SS6[35][21] = 4'h0;
    SS6[36][21] = 4'h0;
    SS6[37][21] = 4'h0;
    SS6[38][21] = 4'h0;
    SS6[39][21] = 4'h0;
    SS6[40][21] = 4'h0;
    SS6[41][21] = 4'h0;
    SS6[42][21] = 4'h0;
    SS6[43][21] = 4'h0;
    SS6[44][21] = 4'h0;
    SS6[45][21] = 4'h0;
    SS6[46][21] = 4'h0;
    SS6[47][21] = 4'h0;
    SS6[0][22] = 4'h0;
    SS6[1][22] = 4'hC;
    SS6[2][22] = 4'hC;
    SS6[3][22] = 4'hC;
    SS6[4][22] = 4'h0;
    SS6[5][22] = 4'h0;
    SS6[6][22] = 4'hC;
    SS6[7][22] = 4'hC;
    SS6[8][22] = 4'hC;
    SS6[9][22] = 4'hC;
    SS6[10][22] = 4'hC;
    SS6[11][22] = 4'hC;
    SS6[12][22] = 4'hC;
    SS6[13][22] = 4'hC;
    SS6[14][22] = 4'hC;
    SS6[15][22] = 4'hC;
    SS6[16][22] = 4'hC;
    SS6[17][22] = 4'hC;
    SS6[18][22] = 4'hD;
    SS6[19][22] = 4'hD;
    SS6[20][22] = 4'hD;
    SS6[21][22] = 4'hC;
    SS6[22][22] = 4'hC;
    SS6[23][22] = 4'hC;
    SS6[24][22] = 4'hC;
    SS6[25][22] = 4'hC;
    SS6[26][22] = 4'hD;
    SS6[27][22] = 4'hC;
    SS6[28][22] = 4'hC;
    SS6[29][22] = 4'hC;
    SS6[30][22] = 4'hD;
    SS6[31][22] = 4'hD;
    SS6[32][22] = 4'hD;
    SS6[33][22] = 4'hD;
    SS6[34][22] = 4'h0;
    SS6[35][22] = 4'h0;
    SS6[36][22] = 4'h0;
    SS6[37][22] = 4'h0;
    SS6[38][22] = 4'h0;
    SS6[39][22] = 4'h0;
    SS6[40][22] = 4'h0;
    SS6[41][22] = 4'h0;
    SS6[42][22] = 4'h0;
    SS6[43][22] = 4'h0;
    SS6[44][22] = 4'h0;
    SS6[45][22] = 4'h0;
    SS6[46][22] = 4'h0;
    SS6[47][22] = 4'h0;
    SS6[0][23] = 4'h0;
    SS6[1][23] = 4'h0;
    SS6[2][23] = 4'hC;
    SS6[3][23] = 4'h0;
    SS6[4][23] = 4'h0;
    SS6[5][23] = 4'h0;
    SS6[6][23] = 4'h0;
    SS6[7][23] = 4'hC;
    SS6[8][23] = 4'hC;
    SS6[9][23] = 4'hC;
    SS6[10][23] = 4'hC;
    SS6[11][23] = 4'hC;
    SS6[12][23] = 4'hC;
    SS6[13][23] = 4'hC;
    SS6[14][23] = 4'hC;
    SS6[15][23] = 4'hC;
    SS6[16][23] = 4'hC;
    SS6[17][23] = 4'hC;
    SS6[18][23] = 4'hC;
    SS6[19][23] = 4'hD;
    SS6[20][23] = 4'hC;
    SS6[21][23] = 4'hC;
    SS6[22][23] = 4'hC;
    SS6[23][23] = 4'hC;
    SS6[24][23] = 4'hC;
    SS6[25][23] = 4'hD;
    SS6[26][23] = 4'hD;
    SS6[27][23] = 4'hD;
    SS6[28][23] = 4'hC;
    SS6[29][23] = 4'hD;
    SS6[30][23] = 4'hD;
    SS6[31][23] = 4'hD;
    SS6[32][23] = 4'hD;
    SS6[33][23] = 4'h0;
    SS6[34][23] = 4'h0;
    SS6[35][23] = 4'h0;
    SS6[36][23] = 4'h0;
    SS6[37][23] = 4'h0;
    SS6[38][23] = 4'h0;
    SS6[39][23] = 4'h0;
    SS6[40][23] = 4'h0;
    SS6[41][23] = 4'h0;
    SS6[42][23] = 4'h0;
    SS6[43][23] = 4'h0;
    SS6[44][23] = 4'h0;
    SS6[45][23] = 4'h0;
    SS6[46][23] = 4'h0;
    SS6[47][23] = 4'h0;
    SS6[0][24] = 4'h0;
    SS6[1][24] = 4'h0;
    SS6[2][24] = 4'h0;
    SS6[3][24] = 4'h0;
    SS6[4][24] = 4'h0;
    SS6[5][24] = 4'h0;
    SS6[6][24] = 4'h0;
    SS6[7][24] = 4'hD;
    SS6[8][24] = 4'hC;
    SS6[9][24] = 4'hC;
    SS6[10][24] = 4'hC;
    SS6[11][24] = 4'hC;
    SS6[12][24] = 4'hC;
    SS6[13][24] = 4'hC;
    SS6[14][24] = 4'hC;
    SS6[15][24] = 4'hC;
    SS6[16][24] = 4'hC;
    SS6[17][24] = 4'hC;
    SS6[18][24] = 4'hC;
    SS6[19][24] = 4'hC;
    SS6[20][24] = 4'hC;
    SS6[21][24] = 4'hC;
    SS6[22][24] = 4'hC;
    SS6[23][24] = 4'hC;
    SS6[24][24] = 4'hD;
    SS6[25][24] = 4'hD;
    SS6[26][24] = 4'hD;
    SS6[27][24] = 4'hD;
    SS6[28][24] = 4'hA;
    SS6[29][24] = 4'hD;
    SS6[30][24] = 4'hD;
    SS6[31][24] = 4'hD;
    SS6[32][24] = 4'hC;
    SS6[33][24] = 4'h0;
    SS6[34][24] = 4'h0;
    SS6[35][24] = 4'h0;
    SS6[36][24] = 4'h0;
    SS6[37][24] = 4'h0;
    SS6[38][24] = 4'h0;
    SS6[39][24] = 4'h0;
    SS6[40][24] = 4'h0;
    SS6[41][24] = 4'h0;
    SS6[42][24] = 4'h0;
    SS6[43][24] = 4'h0;
    SS6[44][24] = 4'h0;
    SS6[45][24] = 4'h0;
    SS6[46][24] = 4'h0;
    SS6[47][24] = 4'h0;
    SS6[0][25] = 4'h0;
    SS6[1][25] = 4'h0;
    SS6[2][25] = 4'h0;
    SS6[3][25] = 4'h0;
    SS6[4][25] = 4'h0;
    SS6[5][25] = 4'h0;
    SS6[6][25] = 4'h0;
    SS6[7][25] = 4'h0;
    SS6[8][25] = 4'hD;
    SS6[9][25] = 4'hC;
    SS6[10][25] = 4'hC;
    SS6[11][25] = 4'hC;
    SS6[12][25] = 4'hC;
    SS6[13][25] = 4'hC;
    SS6[14][25] = 4'hC;
    SS6[15][25] = 4'hC;
    SS6[16][25] = 4'hC;
    SS6[17][25] = 4'hC;
    SS6[18][25] = 4'hC;
    SS6[19][25] = 4'hC;
    SS6[20][25] = 4'hC;
    SS6[21][25] = 4'hC;
    SS6[22][25] = 4'hC;
    SS6[23][25] = 4'hD;
    SS6[24][25] = 4'hD;
    SS6[25][25] = 4'hD;
    SS6[26][25] = 4'hD;
    SS6[27][25] = 4'hA;
    SS6[28][25] = 4'hA;
    SS6[29][25] = 4'hA;
    SS6[30][25] = 4'hD;
    SS6[31][25] = 4'hC;
    SS6[32][25] = 4'hC;
    SS6[33][25] = 4'hC;
    SS6[34][25] = 4'h0;
    SS6[35][25] = 4'h0;
    SS6[36][25] = 4'h0;
    SS6[37][25] = 4'h0;
    SS6[38][25] = 4'h0;
    SS6[39][25] = 4'h0;
    SS6[40][25] = 4'h0;
    SS6[41][25] = 4'h0;
    SS6[42][25] = 4'h0;
    SS6[43][25] = 4'h0;
    SS6[44][25] = 4'h0;
    SS6[45][25] = 4'h0;
    SS6[46][25] = 4'h0;
    SS6[47][25] = 4'h0;
    SS6[0][26] = 4'h0;
    SS6[1][26] = 4'h0;
    SS6[2][26] = 4'h0;
    SS6[3][26] = 4'h0;
    SS6[4][26] = 4'h0;
    SS6[5][26] = 4'h0;
    SS6[6][26] = 4'h0;
    SS6[7][26] = 4'h0;
    SS6[8][26] = 4'h0;
    SS6[9][26] = 4'hE;
    SS6[10][26] = 4'hC;
    SS6[11][26] = 4'hC;
    SS6[12][26] = 4'hC;
    SS6[13][26] = 4'hE;
    SS6[14][26] = 4'hC;
    SS6[15][26] = 4'hC;
    SS6[16][26] = 4'hC;
    SS6[17][26] = 4'hE;
    SS6[18][26] = 4'hC;
    SS6[19][26] = 4'hC;
    SS6[20][26] = 4'hC;
    SS6[21][26] = 4'hC;
    SS6[22][26] = 4'hD;
    SS6[23][26] = 4'hD;
    SS6[24][26] = 4'hD;
    SS6[25][26] = 4'hD;
    SS6[26][26] = 4'hA;
    SS6[27][26] = 4'hA;
    SS6[28][26] = 4'hA;
    SS6[29][26] = 4'hA;
    SS6[30][26] = 4'hC;
    SS6[31][26] = 4'hC;
    SS6[32][26] = 4'hC;
    SS6[33][26] = 4'hC;
    SS6[34][26] = 4'hD;
    SS6[35][26] = 4'h0;
    SS6[36][26] = 4'h0;
    SS6[37][26] = 4'h0;
    SS6[38][26] = 4'h0;
    SS6[39][26] = 4'h0;
    SS6[40][26] = 4'h0;
    SS6[41][26] = 4'h0;
    SS6[42][26] = 4'h0;
    SS6[43][26] = 4'h0;
    SS6[44][26] = 4'h0;
    SS6[45][26] = 4'h0;
    SS6[46][26] = 4'h0;
    SS6[47][26] = 4'h0;
    SS6[0][27] = 4'h0;
    SS6[1][27] = 4'h0;
    SS6[2][27] = 4'h0;
    SS6[3][27] = 4'h0;
    SS6[4][27] = 4'h0;
    SS6[5][27] = 4'h0;
    SS6[6][27] = 4'h0;
    SS6[7][27] = 4'h0;
    SS6[8][27] = 4'hE;
    SS6[9][27] = 4'hE;
    SS6[10][27] = 4'hE;
    SS6[11][27] = 4'hC;
    SS6[12][27] = 4'hE;
    SS6[13][27] = 4'hE;
    SS6[14][27] = 4'hE;
    SS6[15][27] = 4'hC;
    SS6[16][27] = 4'hE;
    SS6[17][27] = 4'hE;
    SS6[18][27] = 4'hE;
    SS6[19][27] = 4'hC;
    SS6[20][27] = 4'hC;
    SS6[21][27] = 4'hC;
    SS6[22][27] = 4'hC;
    SS6[23][27] = 4'hD;
    SS6[24][27] = 4'hD;
    SS6[25][27] = 4'hA;
    SS6[26][27] = 4'hA;
    SS6[27][27] = 4'hA;
    SS6[28][27] = 4'hA;
    SS6[29][27] = 4'hC;
    SS6[30][27] = 4'hC;
    SS6[31][27] = 4'hC;
    SS6[32][27] = 4'hC;
    SS6[33][27] = 4'hD;
    SS6[34][27] = 4'hD;
    SS6[35][27] = 4'hD;
    SS6[36][27] = 4'h0;
    SS6[37][27] = 4'h0;
    SS6[38][27] = 4'h0;
    SS6[39][27] = 4'h0;
    SS6[40][27] = 4'h0;
    SS6[41][27] = 4'h0;
    SS6[42][27] = 4'h0;
    SS6[43][27] = 4'h0;
    SS6[44][27] = 4'h0;
    SS6[45][27] = 4'h0;
    SS6[46][27] = 4'h0;
    SS6[47][27] = 4'h0;
    SS6[0][28] = 4'h0;
    SS6[1][28] = 4'h0;
    SS6[2][28] = 4'h0;
    SS6[3][28] = 4'h0;
    SS6[4][28] = 4'h0;
    SS6[5][28] = 4'h0;
    SS6[6][28] = 4'h0;
    SS6[7][28] = 4'hE;
    SS6[8][28] = 4'hE;
    SS6[9][28] = 4'hE;
    SS6[10][28] = 4'hE;
    SS6[11][28] = 4'hE;
    SS6[12][28] = 4'hE;
    SS6[13][28] = 4'hE;
    SS6[14][28] = 4'hE;
    SS6[15][28] = 4'hD;
    SS6[16][28] = 4'hE;
    SS6[17][28] = 4'hE;
    SS6[18][28] = 4'hE;
    SS6[19][28] = 4'hD;
    SS6[20][28] = 4'hC;
    SS6[21][28] = 4'hC;
    SS6[22][28] = 4'hC;
    SS6[23][28] = 4'hC;
    SS6[24][28] = 4'hA;
    SS6[25][28] = 4'hA;
    SS6[26][28] = 4'hA;
    SS6[27][28] = 4'hA;
    SS6[28][28] = 4'hC;
    SS6[29][28] = 4'hC;
    SS6[30][28] = 4'hC;
    SS6[31][28] = 4'hC;
    SS6[32][28] = 4'hC;
    SS6[33][28] = 4'hD;
    SS6[34][28] = 4'hD;
    SS6[35][28] = 4'hD;
    SS6[36][28] = 4'hD;
    SS6[37][28] = 4'h0;
    SS6[38][28] = 4'h0;
    SS6[39][28] = 4'h0;
    SS6[40][28] = 4'h0;
    SS6[41][28] = 4'h0;
    SS6[42][28] = 4'h0;
    SS6[43][28] = 4'h0;
    SS6[44][28] = 4'h0;
    SS6[45][28] = 4'h0;
    SS6[46][28] = 4'h0;
    SS6[47][28] = 4'h0;
    SS6[0][29] = 4'h0;
    SS6[1][29] = 4'h0;
    SS6[2][29] = 4'h0;
    SS6[3][29] = 4'h0;
    SS6[4][29] = 4'h0;
    SS6[5][29] = 4'h0;
    SS6[6][29] = 4'hE;
    SS6[7][29] = 4'hE;
    SS6[8][29] = 4'hE;
    SS6[9][29] = 4'hE;
    SS6[10][29] = 4'hE;
    SS6[11][29] = 4'hE;
    SS6[12][29] = 4'hE;
    SS6[13][29] = 4'hE;
    SS6[14][29] = 4'hD;
    SS6[15][29] = 4'hD;
    SS6[16][29] = 4'hD;
    SS6[17][29] = 4'hE;
    SS6[18][29] = 4'hD;
    SS6[19][29] = 4'hD;
    SS6[20][29] = 4'hD;
    SS6[21][29] = 4'hC;
    SS6[22][29] = 4'hC;
    SS6[23][29] = 4'hD;
    SS6[24][29] = 4'hD;
    SS6[25][29] = 4'hA;
    SS6[26][29] = 4'hA;
    SS6[27][29] = 4'hC;
    SS6[28][29] = 4'hC;
    SS6[29][29] = 4'hC;
    SS6[30][29] = 4'hC;
    SS6[31][29] = 4'hC;
    SS6[32][29] = 4'hC;
    SS6[33][29] = 4'hC;
    SS6[34][29] = 4'hD;
    SS6[35][29] = 4'hD;
    SS6[36][29] = 4'hD;
    SS6[37][29] = 4'hD;
    SS6[38][29] = 4'h0;
    SS6[39][29] = 4'h0;
    SS6[40][29] = 4'h0;
    SS6[41][29] = 4'h0;
    SS6[42][29] = 4'h0;
    SS6[43][29] = 4'h0;
    SS6[44][29] = 4'h0;
    SS6[45][29] = 4'h0;
    SS6[46][29] = 4'h0;
    SS6[47][29] = 4'h0;
    SS6[0][30] = 4'h0;
    SS6[1][30] = 4'h0;
    SS6[2][30] = 4'h0;
    SS6[3][30] = 4'h0;
    SS6[4][30] = 4'h0;
    SS6[5][30] = 4'hE;
    SS6[6][30] = 4'hE;
    SS6[7][30] = 4'hE;
    SS6[8][30] = 4'hE;
    SS6[9][30] = 4'hE;
    SS6[10][30] = 4'hE;
    SS6[11][30] = 4'hE;
    SS6[12][30] = 4'hE;
    SS6[13][30] = 4'hD;
    SS6[14][30] = 4'hD;
    SS6[15][30] = 4'hD;
    SS6[16][30] = 4'hD;
    SS6[17][30] = 4'hD;
    SS6[18][30] = 4'hD;
    SS6[19][30] = 4'hD;
    SS6[20][30] = 4'hD;
    SS6[21][30] = 4'hD;
    SS6[22][30] = 4'hD;
    SS6[23][30] = 4'hD;
    SS6[24][30] = 4'hD;
    SS6[25][30] = 4'hD;
    SS6[26][30] = 4'hC;
    SS6[27][30] = 4'hC;
    SS6[28][30] = 4'hC;
    SS6[29][30] = 4'hC;
    SS6[30][30] = 4'hC;
    SS6[31][30] = 4'hC;
    SS6[32][30] = 4'hC;
    SS6[33][30] = 4'hC;
    SS6[34][30] = 4'hC;
    SS6[35][30] = 4'hD;
    SS6[36][30] = 4'hD;
    SS6[37][30] = 4'hD;
    SS6[38][30] = 4'hD;
    SS6[39][30] = 4'h0;
    SS6[40][30] = 4'h0;
    SS6[41][30] = 4'h0;
    SS6[42][30] = 4'h0;
    SS6[43][30] = 4'h0;
    SS6[44][30] = 4'h0;
    SS6[45][30] = 4'h0;
    SS6[46][30] = 4'h0;
    SS6[47][30] = 4'h0;
    SS6[0][31] = 4'h0;
    SS6[1][31] = 4'h0;
    SS6[2][31] = 4'h0;
    SS6[3][31] = 4'h0;
    SS6[4][31] = 4'hD;
    SS6[5][31] = 4'hD;
    SS6[6][31] = 4'hE;
    SS6[7][31] = 4'hE;
    SS6[8][31] = 4'hD;
    SS6[9][31] = 4'hD;
    SS6[10][31] = 4'hE;
    SS6[11][31] = 4'hE;
    SS6[12][31] = 4'hD;
    SS6[13][31] = 4'hD;
    SS6[14][31] = 4'hD;
    SS6[15][31] = 4'hD;
    SS6[16][31] = 4'hD;
    SS6[17][31] = 4'hD;
    SS6[18][31] = 4'hD;
    SS6[19][31] = 4'hD;
    SS6[20][31] = 4'hD;
    SS6[21][31] = 4'hD;
    SS6[22][31] = 4'hD;
    SS6[23][31] = 4'hD;
    SS6[24][31] = 4'hD;
    SS6[25][31] = 4'hC;
    SS6[26][31] = 4'hC;
    SS6[27][31] = 4'hC;
    SS6[28][31] = 4'hC;
    SS6[29][31] = 4'hC;
    SS6[30][31] = 4'hC;
    SS6[31][31] = 4'hC;
    SS6[32][31] = 4'hC;
    SS6[33][31] = 4'hC;
    SS6[34][31] = 4'hC;
    SS6[35][31] = 4'hC;
    SS6[36][31] = 4'hD;
    SS6[37][31] = 4'hD;
    SS6[38][31] = 4'hD;
    SS6[39][31] = 4'hD;
    SS6[40][31] = 4'h0;
    SS6[41][31] = 4'h0;
    SS6[42][31] = 4'h0;
    SS6[43][31] = 4'h0;
    SS6[44][31] = 4'h0;
    SS6[45][31] = 4'h0;
    SS6[46][31] = 4'h0;
    SS6[47][31] = 4'h0;
    SS6[0][32] = 4'h0;
    SS6[1][32] = 4'h0;
    SS6[2][32] = 4'h0;
    SS6[3][32] = 4'hD;
    SS6[4][32] = 4'hD;
    SS6[5][32] = 4'hD;
    SS6[6][32] = 4'hD;
    SS6[7][32] = 4'hD;
    SS6[8][32] = 4'hD;
    SS6[9][32] = 4'hD;
    SS6[10][32] = 4'hD;
    SS6[11][32] = 4'hD;
    SS6[12][32] = 4'hD;
    SS6[13][32] = 4'hD;
    SS6[14][32] = 4'hD;
    SS6[15][32] = 4'hD;
    SS6[16][32] = 4'hD;
    SS6[17][32] = 4'hD;
    SS6[18][32] = 4'hD;
    SS6[19][32] = 4'hD;
    SS6[20][32] = 4'hD;
    SS6[21][32] = 4'hD;
    SS6[22][32] = 4'hD;
    SS6[23][32] = 4'hD;
    SS6[24][32] = 4'hC;
    SS6[25][32] = 4'hC;
    SS6[26][32] = 4'hC;
    SS6[27][32] = 4'hC;
    SS6[28][32] = 4'hC;
    SS6[29][32] = 4'hC;
    SS6[30][32] = 4'hC;
    SS6[31][32] = 4'hC;
    SS6[32][32] = 4'hC;
    SS6[33][32] = 4'hC;
    SS6[34][32] = 4'hC;
    SS6[35][32] = 4'hC;
    SS6[36][32] = 4'hC;
    SS6[37][32] = 4'hD;
    SS6[38][32] = 4'hD;
    SS6[39][32] = 4'hD;
    SS6[40][32] = 4'hD;
    SS6[41][32] = 4'h0;
    SS6[42][32] = 4'h0;
    SS6[43][32] = 4'h0;
    SS6[44][32] = 4'h0;
    SS6[45][32] = 4'h0;
    SS6[46][32] = 4'h0;
    SS6[47][32] = 4'h0;
    SS6[0][33] = 4'h0;
    SS6[1][33] = 4'h0;
    SS6[2][33] = 4'hD;
    SS6[3][33] = 4'hD;
    SS6[4][33] = 4'hD;
    SS6[5][33] = 4'hD;
    SS6[6][33] = 4'hD;
    SS6[7][33] = 4'hD;
    SS6[8][33] = 4'hD;
    SS6[9][33] = 4'hD;
    SS6[10][33] = 4'h3;
    SS6[11][33] = 4'h3;
    SS6[12][33] = 4'hD;
    SS6[13][33] = 4'hD;
    SS6[14][33] = 4'hE;
    SS6[15][33] = 4'h0;
    SS6[16][33] = 4'h0;
    SS6[17][33] = 4'hD;
    SS6[18][33] = 4'hD;
    SS6[19][33] = 4'h3;
    SS6[20][33] = 4'h3;
    SS6[21][33] = 4'hD;
    SS6[22][33] = 4'hD;
    SS6[23][33] = 4'h0;
    SS6[24][33] = 4'h0;
    SS6[25][33] = 4'hC;
    SS6[26][33] = 4'hC;
    SS6[27][33] = 4'hD;
    SS6[28][33] = 4'hD;
    SS6[29][33] = 4'hC;
    SS6[30][33] = 4'hC;
    SS6[31][33] = 4'hC;
    SS6[32][33] = 4'hC;
    SS6[33][33] = 4'hC;
    SS6[34][33] = 4'hC;
    SS6[35][33] = 4'hC;
    SS6[36][33] = 4'hC;
    SS6[37][33] = 4'hC;
    SS6[38][33] = 4'hD;
    SS6[39][33] = 4'hD;
    SS6[40][33] = 4'h0;
    SS6[41][33] = 4'h0;
    SS6[42][33] = 4'h0;
    SS6[43][33] = 4'h0;
    SS6[44][33] = 4'h0;
    SS6[45][33] = 4'h0;
    SS6[46][33] = 4'h0;
    SS6[47][33] = 4'h0;
    SS6[0][34] = 4'h0;
    SS6[1][34] = 4'hD;
    SS6[2][34] = 4'hD;
    SS6[3][34] = 4'hD;
    SS6[4][34] = 4'hD;
    SS6[5][34] = 4'hD;
    SS6[6][34] = 4'hD;
    SS6[7][34] = 4'hD;
    SS6[8][34] = 4'hD;
    SS6[9][34] = 4'h3;
    SS6[10][34] = 4'h3;
    SS6[11][34] = 4'h3;
    SS6[12][34] = 4'h3;
    SS6[13][34] = 4'hE;
    SS6[14][34] = 4'h0;
    SS6[15][34] = 4'h0;
    SS6[16][34] = 4'h0;
    SS6[17][34] = 4'h0;
    SS6[18][34] = 4'h3;
    SS6[19][34] = 4'h3;
    SS6[20][34] = 4'h3;
    SS6[21][34] = 4'h3;
    SS6[22][34] = 4'h0;
    SS6[23][34] = 4'h0;
    SS6[24][34] = 4'h0;
    SS6[25][34] = 4'h0;
    SS6[26][34] = 4'hD;
    SS6[27][34] = 4'hD;
    SS6[28][34] = 4'hD;
    SS6[29][34] = 4'hD;
    SS6[30][34] = 4'hC;
    SS6[31][34] = 4'hC;
    SS6[32][34] = 4'hC;
    SS6[33][34] = 4'hC;
    SS6[34][34] = 4'hC;
    SS6[35][34] = 4'hC;
    SS6[36][34] = 4'hC;
    SS6[37][34] = 4'hC;
    SS6[38][34] = 4'hC;
    SS6[39][34] = 4'h0;
    SS6[40][34] = 4'h0;
    SS6[41][34] = 4'h0;
    SS6[42][34] = 4'h0;
    SS6[43][34] = 4'h0;
    SS6[44][34] = 4'h0;
    SS6[45][34] = 4'h0;
    SS6[46][34] = 4'h0;
    SS6[47][34] = 4'h0;
    SS6[0][35] = 4'h0;
    SS6[1][35] = 4'h0;
    SS6[2][35] = 4'hD;
    SS6[3][35] = 4'hD;
    SS6[4][35] = 4'h0;
    SS6[5][35] = 4'h0;
    SS6[6][35] = 4'hD;
    SS6[7][35] = 4'hD;
    SS6[8][35] = 4'h0;
    SS6[9][35] = 4'h0;
    SS6[10][35] = 4'h3;
    SS6[11][35] = 4'h3;
    SS6[12][35] = 4'h2;
    SS6[13][35] = 4'h0;
    SS6[14][35] = 4'h0;
    SS6[15][35] = 4'h0;
    SS6[16][35] = 4'h0;
    SS6[17][35] = 4'h0;
    SS6[18][35] = 4'h2;
    SS6[19][35] = 4'h3;
    SS6[20][35] = 4'h3;
    SS6[21][35] = 4'h0;
    SS6[22][35] = 4'h0;
    SS6[23][35] = 4'h0;
    SS6[24][35] = 4'h0;
    SS6[25][35] = 4'h0;
    SS6[26][35] = 4'h0;
    SS6[27][35] = 4'hD;
    SS6[28][35] = 4'hD;
    SS6[29][35] = 4'hD;
    SS6[30][35] = 4'hD;
    SS6[31][35] = 4'hC;
    SS6[32][35] = 4'hC;
    SS6[33][35] = 4'hC;
    SS6[34][35] = 4'hC;
    SS6[35][35] = 4'hC;
    SS6[36][35] = 4'hC;
    SS6[37][35] = 4'hC;
    SS6[38][35] = 4'hC;
    SS6[39][35] = 4'hC;
    SS6[40][35] = 4'h0;
    SS6[41][35] = 4'h0;
    SS6[42][35] = 4'h0;
    SS6[43][35] = 4'h0;
    SS6[44][35] = 4'h0;
    SS6[45][35] = 4'h0;
    SS6[46][35] = 4'h0;
    SS6[47][35] = 4'h0;
    SS6[0][36] = 4'h0;
    SS6[1][36] = 4'h0;
    SS6[2][36] = 4'h0;
    SS6[3][36] = 4'h0;
    SS6[4][36] = 4'h0;
    SS6[5][36] = 4'h0;
    SS6[6][36] = 4'h0;
    SS6[7][36] = 4'h0;
    SS6[8][36] = 4'h0;
    SS6[9][36] = 4'h0;
    SS6[10][36] = 4'h0;
    SS6[11][36] = 4'h2;
    SS6[12][36] = 4'h0;
    SS6[13][36] = 4'h0;
    SS6[14][36] = 4'h0;
    SS6[15][36] = 4'h0;
    SS6[16][36] = 4'h0;
    SS6[17][36] = 4'h0;
    SS6[18][36] = 4'h0;
    SS6[19][36] = 4'h2;
    SS6[20][36] = 4'h0;
    SS6[21][36] = 4'h0;
    SS6[22][36] = 4'h0;
    SS6[23][36] = 4'h0;
    SS6[24][36] = 4'h0;
    SS6[25][36] = 4'h0;
    SS6[26][36] = 4'h0;
    SS6[27][36] = 4'h0;
    SS6[28][36] = 4'hD;
    SS6[29][36] = 4'hD;
    SS6[30][36] = 4'hD;
    SS6[31][36] = 4'hD;
    SS6[32][36] = 4'hC;
    SS6[33][36] = 4'hC;
    SS6[34][36] = 4'hC;
    SS6[35][36] = 4'hC;
    SS6[36][36] = 4'hC;
    SS6[37][36] = 4'hC;
    SS6[38][36] = 4'hC;
    SS6[39][36] = 4'hC;
    SS6[40][36] = 4'hC;
    SS6[41][36] = 4'h0;
    SS6[42][36] = 4'h0;
    SS6[43][36] = 4'h0;
    SS6[44][36] = 4'h0;
    SS6[45][36] = 4'h0;
    SS6[46][36] = 4'h0;
    SS6[47][36] = 4'h0;
    SS6[0][37] = 4'h0;
    SS6[1][37] = 4'h0;
    SS6[2][37] = 4'h0;
    SS6[3][37] = 4'h0;
    SS6[4][37] = 4'h0;
    SS6[5][37] = 4'h0;
    SS6[6][37] = 4'h0;
    SS6[7][37] = 4'h0;
    SS6[8][37] = 4'h0;
    SS6[9][37] = 4'h0;
    SS6[10][37] = 4'h0;
    SS6[11][37] = 4'h0;
    SS6[12][37] = 4'h0;
    SS6[13][37] = 4'h0;
    SS6[14][37] = 4'h0;
    SS6[15][37] = 4'h0;
    SS6[16][37] = 4'h0;
    SS6[17][37] = 4'h0;
    SS6[18][37] = 4'h0;
    SS6[19][37] = 4'h0;
    SS6[20][37] = 4'h0;
    SS6[21][37] = 4'h0;
    SS6[22][37] = 4'h0;
    SS6[23][37] = 4'h0;
    SS6[24][37] = 4'h0;
    SS6[25][37] = 4'h0;
    SS6[26][37] = 4'h0;
    SS6[27][37] = 4'h0;
    SS6[28][37] = 4'h0;
    SS6[29][37] = 4'hD;
    SS6[30][37] = 4'hD;
    SS6[31][37] = 4'hD;
    SS6[32][37] = 4'hD;
    SS6[33][37] = 4'hC;
    SS6[34][37] = 4'hC;
    SS6[35][37] = 4'hC;
    SS6[36][37] = 4'hC;
    SS6[37][37] = 4'hC;
    SS6[38][37] = 4'hC;
    SS6[39][37] = 4'hC;
    SS6[40][37] = 4'hC;
    SS6[41][37] = 4'hC;
    SS6[42][37] = 4'h0;
    SS6[43][37] = 4'h0;
    SS6[44][37] = 4'h0;
    SS6[45][37] = 4'h0;
    SS6[46][37] = 4'h0;
    SS6[47][37] = 4'h0;
    SS6[0][38] = 4'h0;
    SS6[1][38] = 4'h0;
    SS6[2][38] = 4'h0;
    SS6[3][38] = 4'h0;
    SS6[4][38] = 4'h0;
    SS6[5][38] = 4'h0;
    SS6[6][38] = 4'h0;
    SS6[7][38] = 4'h0;
    SS6[8][38] = 4'h0;
    SS6[9][38] = 4'h0;
    SS6[10][38] = 4'h0;
    SS6[11][38] = 4'h0;
    SS6[12][38] = 4'h0;
    SS6[13][38] = 4'h0;
    SS6[14][38] = 4'h0;
    SS6[15][38] = 4'h0;
    SS6[16][38] = 4'h0;
    SS6[17][38] = 4'h0;
    SS6[18][38] = 4'h0;
    SS6[19][38] = 4'h0;
    SS6[20][38] = 4'h0;
    SS6[21][38] = 4'h0;
    SS6[22][38] = 4'h0;
    SS6[23][38] = 4'h0;
    SS6[24][38] = 4'h0;
    SS6[25][38] = 4'h0;
    SS6[26][38] = 4'h0;
    SS6[27][38] = 4'h0;
    SS6[28][38] = 4'h0;
    SS6[29][38] = 4'h0;
    SS6[30][38] = 4'hD;
    SS6[31][38] = 4'hD;
    SS6[32][38] = 4'hD;
    SS6[33][38] = 4'hD;
    SS6[34][38] = 4'hC;
    SS6[35][38] = 4'hC;
    SS6[36][38] = 4'hC;
    SS6[37][38] = 4'hC;
    SS6[38][38] = 4'hC;
    SS6[39][38] = 4'hC;
    SS6[40][38] = 4'hC;
    SS6[41][38] = 4'hC;
    SS6[42][38] = 4'hC;
    SS6[43][38] = 4'h0;
    SS6[44][38] = 4'h0;
    SS6[45][38] = 4'h0;
    SS6[46][38] = 4'h0;
    SS6[47][38] = 4'h0;
    SS6[0][39] = 4'h0;
    SS6[1][39] = 4'h0;
    SS6[2][39] = 4'h0;
    SS6[3][39] = 4'h0;
    SS6[4][39] = 4'h0;
    SS6[5][39] = 4'h0;
    SS6[6][39] = 4'h0;
    SS6[7][39] = 4'h0;
    SS6[8][39] = 4'h0;
    SS6[9][39] = 4'h0;
    SS6[10][39] = 4'h0;
    SS6[11][39] = 4'h0;
    SS6[12][39] = 4'h0;
    SS6[13][39] = 4'h0;
    SS6[14][39] = 4'h0;
    SS6[15][39] = 4'h0;
    SS6[16][39] = 4'h0;
    SS6[17][39] = 4'h0;
    SS6[18][39] = 4'h0;
    SS6[19][39] = 4'h0;
    SS6[20][39] = 4'h0;
    SS6[21][39] = 4'h0;
    SS6[22][39] = 4'h0;
    SS6[23][39] = 4'h0;
    SS6[24][39] = 4'h0;
    SS6[25][39] = 4'h0;
    SS6[26][39] = 4'h0;
    SS6[27][39] = 4'h0;
    SS6[28][39] = 4'h0;
    SS6[29][39] = 4'h0;
    SS6[30][39] = 4'h0;
    SS6[31][39] = 4'hD;
    SS6[32][39] = 4'hD;
    SS6[33][39] = 4'hD;
    SS6[34][39] = 4'h0;
    SS6[35][39] = 4'hC;
    SS6[36][39] = 4'hC;
    SS6[37][39] = 4'hC;
    SS6[38][39] = 4'hC;
    SS6[39][39] = 4'hC;
    SS6[40][39] = 4'hC;
    SS6[41][39] = 4'hC;
    SS6[42][39] = 4'h0;
    SS6[43][39] = 4'h0;
    SS6[44][39] = 4'h0;
    SS6[45][39] = 4'h0;
    SS6[46][39] = 4'h0;
    SS6[47][39] = 4'h0;
    SS6[0][40] = 4'h0;
    SS6[1][40] = 4'h0;
    SS6[2][40] = 4'h0;
    SS6[3][40] = 4'h0;
    SS6[4][40] = 4'h0;
    SS6[5][40] = 4'h0;
    SS6[6][40] = 4'h0;
    SS6[7][40] = 4'h0;
    SS6[8][40] = 4'h0;
    SS6[9][40] = 4'h0;
    SS6[10][40] = 4'h0;
    SS6[11][40] = 4'h0;
    SS6[12][40] = 4'h0;
    SS6[13][40] = 4'h0;
    SS6[14][40] = 4'h0;
    SS6[15][40] = 4'h0;
    SS6[16][40] = 4'h0;
    SS6[17][40] = 4'h0;
    SS6[18][40] = 4'h0;
    SS6[19][40] = 4'h0;
    SS6[20][40] = 4'h0;
    SS6[21][40] = 4'h0;
    SS6[22][40] = 4'h0;
    SS6[23][40] = 4'h0;
    SS6[24][40] = 4'h0;
    SS6[25][40] = 4'h0;
    SS6[26][40] = 4'h0;
    SS6[27][40] = 4'h0;
    SS6[28][40] = 4'h0;
    SS6[29][40] = 4'h0;
    SS6[30][40] = 4'h0;
    SS6[31][40] = 4'h0;
    SS6[32][40] = 4'hD;
    SS6[33][40] = 4'h0;
    SS6[34][40] = 4'h0;
    SS6[35][40] = 4'h0;
    SS6[36][40] = 4'hC;
    SS6[37][40] = 4'hC;
    SS6[38][40] = 4'hC;
    SS6[39][40] = 4'hC;
    SS6[40][40] = 4'hC;
    SS6[41][40] = 4'h0;
    SS6[42][40] = 4'h0;
    SS6[43][40] = 4'h0;
    SS6[44][40] = 4'h0;
    SS6[45][40] = 4'h0;
    SS6[46][40] = 4'h0;
    SS6[47][40] = 4'h0;
    SS6[0][41] = 4'h0;
    SS6[1][41] = 4'h0;
    SS6[2][41] = 4'h0;
    SS6[3][41] = 4'h0;
    SS6[4][41] = 4'h0;
    SS6[5][41] = 4'h0;
    SS6[6][41] = 4'h0;
    SS6[7][41] = 4'h0;
    SS6[8][41] = 4'h0;
    SS6[9][41] = 4'h0;
    SS6[10][41] = 4'h0;
    SS6[11][41] = 4'h0;
    SS6[12][41] = 4'h0;
    SS6[13][41] = 4'h0;
    SS6[14][41] = 4'h0;
    SS6[15][41] = 4'h0;
    SS6[16][41] = 4'h0;
    SS6[17][41] = 4'h0;
    SS6[18][41] = 4'h0;
    SS6[19][41] = 4'h0;
    SS6[20][41] = 4'h0;
    SS6[21][41] = 4'h0;
    SS6[22][41] = 4'h0;
    SS6[23][41] = 4'h0;
    SS6[24][41] = 4'h0;
    SS6[25][41] = 4'h0;
    SS6[26][41] = 4'h0;
    SS6[27][41] = 4'h0;
    SS6[28][41] = 4'h0;
    SS6[29][41] = 4'h0;
    SS6[30][41] = 4'h0;
    SS6[31][41] = 4'h0;
    SS6[32][41] = 4'h0;
    SS6[33][41] = 4'h0;
    SS6[34][41] = 4'h0;
    SS6[35][41] = 4'h0;
    SS6[36][41] = 4'h0;
    SS6[37][41] = 4'hC;
    SS6[38][41] = 4'hC;
    SS6[39][41] = 4'hC;
    SS6[40][41] = 4'h0;
    SS6[41][41] = 4'h0;
    SS6[42][41] = 4'h0;
    SS6[43][41] = 4'h0;
    SS6[44][41] = 4'h0;
    SS6[45][41] = 4'h0;
    SS6[46][41] = 4'h0;
    SS6[47][41] = 4'h0;
    SS6[0][42] = 4'h0;
    SS6[1][42] = 4'h0;
    SS6[2][42] = 4'h0;
    SS6[3][42] = 4'h0;
    SS6[4][42] = 4'h0;
    SS6[5][42] = 4'h0;
    SS6[6][42] = 4'h0;
    SS6[7][42] = 4'h0;
    SS6[8][42] = 4'h0;
    SS6[9][42] = 4'h0;
    SS6[10][42] = 4'h0;
    SS6[11][42] = 4'h0;
    SS6[12][42] = 4'h0;
    SS6[13][42] = 4'h0;
    SS6[14][42] = 4'h0;
    SS6[15][42] = 4'h0;
    SS6[16][42] = 4'h0;
    SS6[17][42] = 4'h0;
    SS6[18][42] = 4'h0;
    SS6[19][42] = 4'h0;
    SS6[20][42] = 4'h0;
    SS6[21][42] = 4'h0;
    SS6[22][42] = 4'h0;
    SS6[23][42] = 4'h0;
    SS6[24][42] = 4'h0;
    SS6[25][42] = 4'h0;
    SS6[26][42] = 4'h0;
    SS6[27][42] = 4'h0;
    SS6[28][42] = 4'h0;
    SS6[29][42] = 4'h0;
    SS6[30][42] = 4'h0;
    SS6[31][42] = 4'h0;
    SS6[32][42] = 4'h0;
    SS6[33][42] = 4'h0;
    SS6[34][42] = 4'h0;
    SS6[35][42] = 4'h0;
    SS6[36][42] = 4'h0;
    SS6[37][42] = 4'h0;
    SS6[38][42] = 4'hC;
    SS6[39][42] = 4'h0;
    SS6[40][42] = 4'h0;
    SS6[41][42] = 4'h0;
    SS6[42][42] = 4'h0;
    SS6[43][42] = 4'h0;
    SS6[44][42] = 4'h0;
    SS6[45][42] = 4'h0;
    SS6[46][42] = 4'h0;
    SS6[47][42] = 4'h0;
    SS6[0][43] = 4'h0;
    SS6[1][43] = 4'h0;
    SS6[2][43] = 4'h0;
    SS6[3][43] = 4'h0;
    SS6[4][43] = 4'h0;
    SS6[5][43] = 4'h0;
    SS6[6][43] = 4'h0;
    SS6[7][43] = 4'h0;
    SS6[8][43] = 4'h0;
    SS6[9][43] = 4'h0;
    SS6[10][43] = 4'h0;
    SS6[11][43] = 4'h0;
    SS6[12][43] = 4'h0;
    SS6[13][43] = 4'h0;
    SS6[14][43] = 4'h0;
    SS6[15][43] = 4'h0;
    SS6[16][43] = 4'h0;
    SS6[17][43] = 4'h0;
    SS6[18][43] = 4'h0;
    SS6[19][43] = 4'h0;
    SS6[20][43] = 4'h0;
    SS6[21][43] = 4'h0;
    SS6[22][43] = 4'h0;
    SS6[23][43] = 4'h0;
    SS6[24][43] = 4'h0;
    SS6[25][43] = 4'h0;
    SS6[26][43] = 4'h0;
    SS6[27][43] = 4'h0;
    SS6[28][43] = 4'h0;
    SS6[29][43] = 4'h0;
    SS6[30][43] = 4'h0;
    SS6[31][43] = 4'h0;
    SS6[32][43] = 4'h0;
    SS6[33][43] = 4'h0;
    SS6[34][43] = 4'h0;
    SS6[35][43] = 4'h0;
    SS6[36][43] = 4'h0;
    SS6[37][43] = 4'h0;
    SS6[38][43] = 4'h0;
    SS6[39][43] = 4'h0;
    SS6[40][43] = 4'h0;
    SS6[41][43] = 4'h0;
    SS6[42][43] = 4'h0;
    SS6[43][43] = 4'h0;
    SS6[44][43] = 4'h0;
    SS6[45][43] = 4'h0;
    SS6[46][43] = 4'h0;
    SS6[47][43] = 4'h0;
    SS6[0][44] = 4'h0;
    SS6[1][44] = 4'h0;
    SS6[2][44] = 4'h0;
    SS6[3][44] = 4'h0;
    SS6[4][44] = 4'h0;
    SS6[5][44] = 4'h0;
    SS6[6][44] = 4'h0;
    SS6[7][44] = 4'h0;
    SS6[8][44] = 4'h0;
    SS6[9][44] = 4'h0;
    SS6[10][44] = 4'h0;
    SS6[11][44] = 4'h0;
    SS6[12][44] = 4'h0;
    SS6[13][44] = 4'h0;
    SS6[14][44] = 4'h0;
    SS6[15][44] = 4'h0;
    SS6[16][44] = 4'h0;
    SS6[17][44] = 4'h0;
    SS6[18][44] = 4'h0;
    SS6[19][44] = 4'h0;
    SS6[20][44] = 4'h0;
    SS6[21][44] = 4'h0;
    SS6[22][44] = 4'h0;
    SS6[23][44] = 4'h0;
    SS6[24][44] = 4'h0;
    SS6[25][44] = 4'h0;
    SS6[26][44] = 4'h0;
    SS6[27][44] = 4'h0;
    SS6[28][44] = 4'h0;
    SS6[29][44] = 4'h0;
    SS6[30][44] = 4'h0;
    SS6[31][44] = 4'h0;
    SS6[32][44] = 4'h0;
    SS6[33][44] = 4'h0;
    SS6[34][44] = 4'h0;
    SS6[35][44] = 4'h0;
    SS6[36][44] = 4'h0;
    SS6[37][44] = 4'h0;
    SS6[38][44] = 4'h0;
    SS6[39][44] = 4'h0;
    SS6[40][44] = 4'h0;
    SS6[41][44] = 4'h0;
    SS6[42][44] = 4'h0;
    SS6[43][44] = 4'h0;
    SS6[44][44] = 4'h0;
    SS6[45][44] = 4'h0;
    SS6[46][44] = 4'h0;
    SS6[47][44] = 4'h0;
    SS6[0][45] = 4'h0;
    SS6[1][45] = 4'h0;
    SS6[2][45] = 4'h0;
    SS6[3][45] = 4'h0;
    SS6[4][45] = 4'h0;
    SS6[5][45] = 4'h0;
    SS6[6][45] = 4'h0;
    SS6[7][45] = 4'h0;
    SS6[8][45] = 4'h0;
    SS6[9][45] = 4'h0;
    SS6[10][45] = 4'h0;
    SS6[11][45] = 4'h0;
    SS6[12][45] = 4'h0;
    SS6[13][45] = 4'h0;
    SS6[14][45] = 4'h0;
    SS6[15][45] = 4'h0;
    SS6[16][45] = 4'h0;
    SS6[17][45] = 4'h0;
    SS6[18][45] = 4'h0;
    SS6[19][45] = 4'h0;
    SS6[20][45] = 4'h0;
    SS6[21][45] = 4'h0;
    SS6[22][45] = 4'h0;
    SS6[23][45] = 4'h0;
    SS6[24][45] = 4'h0;
    SS6[25][45] = 4'h0;
    SS6[26][45] = 4'h0;
    SS6[27][45] = 4'h0;
    SS6[28][45] = 4'h0;
    SS6[29][45] = 4'h0;
    SS6[30][45] = 4'h0;
    SS6[31][45] = 4'h0;
    SS6[32][45] = 4'h0;
    SS6[33][45] = 4'h0;
    SS6[34][45] = 4'h0;
    SS6[35][45] = 4'h0;
    SS6[36][45] = 4'h0;
    SS6[37][45] = 4'h0;
    SS6[38][45] = 4'h0;
    SS6[39][45] = 4'h0;
    SS6[40][45] = 4'h0;
    SS6[41][45] = 4'h0;
    SS6[42][45] = 4'h0;
    SS6[43][45] = 4'h0;
    SS6[44][45] = 4'h0;
    SS6[45][45] = 4'h0;
    SS6[46][45] = 4'h0;
    SS6[47][45] = 4'h0;
    SS6[0][46] = 4'h0;
    SS6[1][46] = 4'h0;
    SS6[2][46] = 4'h0;
    SS6[3][46] = 4'h0;
    SS6[4][46] = 4'h0;
    SS6[5][46] = 4'h0;
    SS6[6][46] = 4'h0;
    SS6[7][46] = 4'h0;
    SS6[8][46] = 4'h0;
    SS6[9][46] = 4'h0;
    SS6[10][46] = 4'h0;
    SS6[11][46] = 4'h0;
    SS6[12][46] = 4'h0;
    SS6[13][46] = 4'h0;
    SS6[14][46] = 4'h0;
    SS6[15][46] = 4'h0;
    SS6[16][46] = 4'h0;
    SS6[17][46] = 4'h0;
    SS6[18][46] = 4'h0;
    SS6[19][46] = 4'h0;
    SS6[20][46] = 4'h0;
    SS6[21][46] = 4'h0;
    SS6[22][46] = 4'h0;
    SS6[23][46] = 4'h0;
    SS6[24][46] = 4'h0;
    SS6[25][46] = 4'h0;
    SS6[26][46] = 4'h0;
    SS6[27][46] = 4'h0;
    SS6[28][46] = 4'h0;
    SS6[29][46] = 4'h0;
    SS6[30][46] = 4'h0;
    SS6[31][46] = 4'h0;
    SS6[32][46] = 4'h0;
    SS6[33][46] = 4'h0;
    SS6[34][46] = 4'h0;
    SS6[35][46] = 4'h0;
    SS6[36][46] = 4'h0;
    SS6[37][46] = 4'h0;
    SS6[38][46] = 4'h0;
    SS6[39][46] = 4'h0;
    SS6[40][46] = 4'h0;
    SS6[41][46] = 4'h0;
    SS6[42][46] = 4'h0;
    SS6[43][46] = 4'h0;
    SS6[44][46] = 4'h0;
    SS6[45][46] = 4'h0;
    SS6[46][46] = 4'h0;
    SS6[47][46] = 4'h0;
    SS6[0][47] = 4'h0;
    SS6[1][47] = 4'h0;
    SS6[2][47] = 4'h0;
    SS6[3][47] = 4'h0;
    SS6[4][47] = 4'h0;
    SS6[5][47] = 4'h0;
    SS6[6][47] = 4'h0;
    SS6[7][47] = 4'h0;
    SS6[8][47] = 4'h0;
    SS6[9][47] = 4'h0;
    SS6[10][47] = 4'h0;
    SS6[11][47] = 4'h0;
    SS6[12][47] = 4'h0;
    SS6[13][47] = 4'h0;
    SS6[14][47] = 4'h0;
    SS6[15][47] = 4'h0;
    SS6[16][47] = 4'h0;
    SS6[17][47] = 4'h0;
    SS6[18][47] = 4'h0;
    SS6[19][47] = 4'h0;
    SS6[20][47] = 4'h0;
    SS6[21][47] = 4'h0;
    SS6[22][47] = 4'h0;
    SS6[23][47] = 4'h0;
    SS6[24][47] = 4'h0;
    SS6[25][47] = 4'h0;
    SS6[26][47] = 4'h0;
    SS6[27][47] = 4'h0;
    SS6[28][47] = 4'h0;
    SS6[29][47] = 4'h0;
    SS6[30][47] = 4'h0;
    SS6[31][47] = 4'h0;
    SS6[32][47] = 4'h0;
    SS6[33][47] = 4'h0;
    SS6[34][47] = 4'h0;
    SS6[35][47] = 4'h0;
    SS6[36][47] = 4'h0;
    SS6[37][47] = 4'h0;
    SS6[38][47] = 4'h0;
    SS6[39][47] = 4'h0;
    SS6[40][47] = 4'h0;
    SS6[41][47] = 4'h0;
    SS6[42][47] = 4'h0;
    SS6[43][47] = 4'h0;
    SS6[44][47] = 4'h0;
    SS6[45][47] = 4'h0;
    SS6[46][47] = 4'h0;
    SS6[47][47] = 4'h0;
 
//SS 7
    SS7[0][0] = 4'h0;
    SS7[1][0] = 4'h0;
    SS7[2][0] = 4'h0;
    SS7[3][0] = 4'h0;
    SS7[4][0] = 4'h0;
    SS7[5][0] = 4'h0;
    SS7[6][0] = 4'h0;
    SS7[7][0] = 4'h0;
    SS7[8][0] = 4'h0;
    SS7[9][0] = 4'h0;
    SS7[10][0] = 4'h0;
    SS7[11][0] = 4'h0;
    SS7[12][0] = 4'h0;
    SS7[13][0] = 4'h0;
    SS7[14][0] = 4'h0;
    SS7[15][0] = 4'h0;
    SS7[16][0] = 4'h0;
    SS7[17][0] = 4'h0;
    SS7[18][0] = 4'h0;
    SS7[19][0] = 4'h0;
    SS7[20][0] = 4'h0;
    SS7[21][0] = 4'h0;
    SS7[22][0] = 4'h0;
    SS7[23][0] = 4'h0;
    SS7[24][0] = 4'h0;
    SS7[25][0] = 4'h0;
    SS7[26][0] = 4'h0;
    SS7[27][0] = 4'hC;
    SS7[28][0] = 4'hC;
    SS7[29][0] = 4'hC;
    SS7[30][0] = 4'h0;
    SS7[31][0] = 4'h0;
    SS7[32][0] = 4'h0;
    SS7[33][0] = 4'h0;
    SS7[34][0] = 4'h0;
    SS7[35][0] = 4'h0;
    SS7[36][0] = 4'h0;
    SS7[37][0] = 4'h0;
    SS7[38][0] = 4'h0;
    SS7[39][0] = 4'h0;
    SS7[40][0] = 4'h0;
    SS7[41][0] = 4'h0;
    SS7[42][0] = 4'h0;
    SS7[43][0] = 4'h0;
    SS7[44][0] = 4'h0;
    SS7[45][0] = 4'h0;
    SS7[46][0] = 4'h0;
    SS7[47][0] = 4'h0;
    SS7[0][1] = 4'h0;
    SS7[1][1] = 4'h0;
    SS7[2][1] = 4'h0;
    SS7[3][1] = 4'h0;
    SS7[4][1] = 4'h0;
    SS7[5][1] = 4'h0;
    SS7[6][1] = 4'h0;
    SS7[7][1] = 4'h0;
    SS7[8][1] = 4'h0;
    SS7[9][1] = 4'h0;
    SS7[10][1] = 4'h0;
    SS7[11][1] = 4'h0;
    SS7[12][1] = 4'h0;
    SS7[13][1] = 4'h0;
    SS7[14][1] = 4'h0;
    SS7[15][1] = 4'h0;
    SS7[16][1] = 4'h0;
    SS7[17][1] = 4'h0;
    SS7[18][1] = 4'h0;
    SS7[19][1] = 4'h0;
    SS7[20][1] = 4'h0;
    SS7[21][1] = 4'h0;
    SS7[22][1] = 4'h0;
    SS7[23][1] = 4'h0;
    SS7[24][1] = 4'hD;
    SS7[25][1] = 4'hD;
    SS7[26][1] = 4'hD;
    SS7[27][1] = 4'hD;
    SS7[28][1] = 4'hC;
    SS7[29][1] = 4'hC;
    SS7[30][1] = 4'hC;
    SS7[31][1] = 4'h0;
    SS7[32][1] = 4'h0;
    SS7[33][1] = 4'h0;
    SS7[34][1] = 4'h0;
    SS7[35][1] = 4'h0;
    SS7[36][1] = 4'h0;
    SS7[37][1] = 4'h0;
    SS7[38][1] = 4'h0;
    SS7[39][1] = 4'h0;
    SS7[40][1] = 4'h0;
    SS7[41][1] = 4'h0;
    SS7[42][1] = 4'h0;
    SS7[43][1] = 4'h0;
    SS7[44][1] = 4'h0;
    SS7[45][1] = 4'h0;
    SS7[46][1] = 4'h0;
    SS7[47][1] = 4'h0;
    SS7[0][2] = 4'h0;
    SS7[1][2] = 4'h0;
    SS7[2][2] = 4'h0;
    SS7[3][2] = 4'h0;
    SS7[4][2] = 4'h0;
    SS7[5][2] = 4'h0;
    SS7[6][2] = 4'h0;
    SS7[7][2] = 4'h0;
    SS7[8][2] = 4'h0;
    SS7[9][2] = 4'h0;
    SS7[10][2] = 4'h0;
    SS7[11][2] = 4'h0;
    SS7[12][2] = 4'h0;
    SS7[13][2] = 4'h0;
    SS7[14][2] = 4'h0;
    SS7[15][2] = 4'h0;
    SS7[16][2] = 4'h0;
    SS7[17][2] = 4'h0;
    SS7[18][2] = 4'h0;
    SS7[19][2] = 4'h0;
    SS7[20][2] = 4'h0;
    SS7[21][2] = 4'h0;
    SS7[22][2] = 4'h0;
    SS7[23][2] = 4'h0;
    SS7[24][2] = 4'h0;
    SS7[25][2] = 4'hD;
    SS7[26][2] = 4'hD;
    SS7[27][2] = 4'hD;
    SS7[28][2] = 4'hC;
    SS7[29][2] = 4'hC;
    SS7[30][2] = 4'hC;
    SS7[31][2] = 4'h0;
    SS7[32][2] = 4'h0;
    SS7[33][2] = 4'h0;
    SS7[34][2] = 4'h0;
    SS7[35][2] = 4'h0;
    SS7[36][2] = 4'h0;
    SS7[37][2] = 4'h0;
    SS7[38][2] = 4'h0;
    SS7[39][2] = 4'h0;
    SS7[40][2] = 4'h0;
    SS7[41][2] = 4'h0;
    SS7[42][2] = 4'h0;
    SS7[43][2] = 4'h0;
    SS7[44][2] = 4'h0;
    SS7[45][2] = 4'h0;
    SS7[46][2] = 4'h0;
    SS7[47][2] = 4'h0;
    SS7[0][3] = 4'h0;
    SS7[1][3] = 4'h0;
    SS7[2][3] = 4'h0;
    SS7[3][3] = 4'h0;
    SS7[4][3] = 4'h0;
    SS7[5][3] = 4'h0;
    SS7[6][3] = 4'h0;
    SS7[7][3] = 4'h0;
    SS7[8][3] = 4'h0;
    SS7[9][3] = 4'h0;
    SS7[10][3] = 4'h0;
    SS7[11][3] = 4'h0;
    SS7[12][3] = 4'h0;
    SS7[13][3] = 4'h0;
    SS7[14][3] = 4'h0;
    SS7[15][3] = 4'h0;
    SS7[16][3] = 4'h0;
    SS7[17][3] = 4'h0;
    SS7[18][3] = 4'h0;
    SS7[19][3] = 4'h0;
    SS7[20][3] = 4'h0;
    SS7[21][3] = 4'h0;
    SS7[22][3] = 4'h0;
    SS7[23][3] = 4'h0;
    SS7[24][3] = 4'h0;
    SS7[25][3] = 4'hD;
    SS7[26][3] = 4'hD;
    SS7[27][3] = 4'hC;
    SS7[28][3] = 4'hC;
    SS7[29][3] = 4'hC;
    SS7[30][3] = 4'hC;
    SS7[31][3] = 4'hC;
    SS7[32][3] = 4'h0;
    SS7[33][3] = 4'h0;
    SS7[34][3] = 4'h0;
    SS7[35][3] = 4'h0;
    SS7[36][3] = 4'h0;
    SS7[37][3] = 4'h0;
    SS7[38][3] = 4'h0;
    SS7[39][3] = 4'h0;
    SS7[40][3] = 4'h0;
    SS7[41][3] = 4'h0;
    SS7[42][3] = 4'h0;
    SS7[43][3] = 4'h0;
    SS7[44][3] = 4'h0;
    SS7[45][3] = 4'h0;
    SS7[46][3] = 4'h0;
    SS7[47][3] = 4'h0;
    SS7[0][4] = 4'h0;
    SS7[1][4] = 4'h0;
    SS7[2][4] = 4'h0;
    SS7[3][4] = 4'h0;
    SS7[4][4] = 4'h0;
    SS7[5][4] = 4'h0;
    SS7[6][4] = 4'h0;
    SS7[7][4] = 4'h0;
    SS7[8][4] = 4'h0;
    SS7[9][4] = 4'h0;
    SS7[10][4] = 4'h0;
    SS7[11][4] = 4'h0;
    SS7[12][4] = 4'h0;
    SS7[13][4] = 4'h0;
    SS7[14][4] = 4'h0;
    SS7[15][4] = 4'h0;
    SS7[16][4] = 4'h0;
    SS7[17][4] = 4'h0;
    SS7[18][4] = 4'h0;
    SS7[19][4] = 4'h0;
    SS7[20][4] = 4'h0;
    SS7[21][4] = 4'h0;
    SS7[22][4] = 4'h0;
    SS7[23][4] = 4'h0;
    SS7[24][4] = 4'h0;
    SS7[25][4] = 4'hE;
    SS7[26][4] = 4'hC;
    SS7[27][4] = 4'hC;
    SS7[28][4] = 4'hC;
    SS7[29][4] = 4'hC;
    SS7[30][4] = 4'hC;
    SS7[31][4] = 4'hC;
    SS7[32][4] = 4'h0;
    SS7[33][4] = 4'h0;
    SS7[34][4] = 4'h0;
    SS7[35][4] = 4'h0;
    SS7[36][4] = 4'h0;
    SS7[37][4] = 4'h0;
    SS7[38][4] = 4'h0;
    SS7[39][4] = 4'h0;
    SS7[40][4] = 4'h0;
    SS7[41][4] = 4'h0;
    SS7[42][4] = 4'h0;
    SS7[43][4] = 4'h0;
    SS7[44][4] = 4'h0;
    SS7[45][4] = 4'h0;
    SS7[46][4] = 4'h0;
    SS7[47][4] = 4'h0;
    SS7[0][5] = 4'h0;
    SS7[1][5] = 4'h0;
    SS7[2][5] = 4'h0;
    SS7[3][5] = 4'h0;
    SS7[4][5] = 4'h0;
    SS7[5][5] = 4'h0;
    SS7[6][5] = 4'h0;
    SS7[7][5] = 4'h0;
    SS7[8][5] = 4'h0;
    SS7[9][5] = 4'h0;
    SS7[10][5] = 4'h0;
    SS7[11][5] = 4'h0;
    SS7[12][5] = 4'h0;
    SS7[13][5] = 4'h0;
    SS7[14][5] = 4'h0;
    SS7[15][5] = 4'h0;
    SS7[16][5] = 4'h0;
    SS7[17][5] = 4'h0;
    SS7[18][5] = 4'h0;
    SS7[19][5] = 4'h0;
    SS7[20][5] = 4'h0;
    SS7[21][5] = 4'h0;
    SS7[22][5] = 4'h0;
    SS7[23][5] = 4'hE;
    SS7[24][5] = 4'hE;
    SS7[25][5] = 4'hE;
    SS7[26][5] = 4'hC;
    SS7[27][5] = 4'hC;
    SS7[28][5] = 4'hC;
    SS7[29][5] = 4'hC;
    SS7[30][5] = 4'h0;
    SS7[31][5] = 4'h0;
    SS7[32][5] = 4'h0;
    SS7[33][5] = 4'h0;
    SS7[34][5] = 4'h0;
    SS7[35][5] = 4'h0;
    SS7[36][5] = 4'h0;
    SS7[37][5] = 4'h0;
    SS7[38][5] = 4'h0;
    SS7[39][5] = 4'h0;
    SS7[40][5] = 4'h0;
    SS7[41][5] = 4'h0;
    SS7[42][5] = 4'h0;
    SS7[43][5] = 4'h0;
    SS7[44][5] = 4'h0;
    SS7[45][5] = 4'h0;
    SS7[46][5] = 4'h0;
    SS7[47][5] = 4'h0;
    SS7[0][6] = 4'h0;
    SS7[1][6] = 4'h0;
    SS7[2][6] = 4'h0;
    SS7[3][6] = 4'h0;
    SS7[4][6] = 4'h0;
    SS7[5][6] = 4'h0;
    SS7[6][6] = 4'h0;
    SS7[7][6] = 4'h0;
    SS7[8][6] = 4'h0;
    SS7[9][6] = 4'h0;
    SS7[10][6] = 4'h0;
    SS7[11][6] = 4'h0;
    SS7[12][6] = 4'h0;
    SS7[13][6] = 4'h0;
    SS7[14][6] = 4'h0;
    SS7[15][6] = 4'h0;
    SS7[16][6] = 4'h0;
    SS7[17][6] = 4'h0;
    SS7[18][6] = 4'h0;
    SS7[19][6] = 4'h0;
    SS7[20][6] = 4'h0;
    SS7[21][6] = 4'h0;
    SS7[22][6] = 4'h0;
    SS7[23][6] = 4'hE;
    SS7[24][6] = 4'hE;
    SS7[25][6] = 4'hE;
    SS7[26][6] = 4'hC;
    SS7[27][6] = 4'hC;
    SS7[28][6] = 4'hC;
    SS7[29][6] = 4'hC;
    SS7[30][6] = 4'h0;
    SS7[31][6] = 4'h0;
    SS7[32][6] = 4'h0;
    SS7[33][6] = 4'h0;
    SS7[34][6] = 4'h0;
    SS7[35][6] = 4'h0;
    SS7[36][6] = 4'h0;
    SS7[37][6] = 4'h0;
    SS7[38][6] = 4'h0;
    SS7[39][6] = 4'h0;
    SS7[40][6] = 4'h0;
    SS7[41][6] = 4'h0;
    SS7[42][6] = 4'h0;
    SS7[43][6] = 4'h0;
    SS7[44][6] = 4'h0;
    SS7[45][6] = 4'h0;
    SS7[46][6] = 4'h0;
    SS7[47][6] = 4'h0;
    SS7[0][7] = 4'h0;
    SS7[1][7] = 4'h0;
    SS7[2][7] = 4'hD;
    SS7[3][7] = 4'hD;
    SS7[4][7] = 4'h0;
    SS7[5][7] = 4'h0;
    SS7[6][7] = 4'h0;
    SS7[7][7] = 4'h0;
    SS7[8][7] = 4'h0;
    SS7[9][7] = 4'h0;
    SS7[10][7] = 4'h0;
    SS7[11][7] = 4'h0;
    SS7[12][7] = 4'h0;
    SS7[13][7] = 4'h0;
    SS7[14][7] = 4'h0;
    SS7[15][7] = 4'h0;
    SS7[16][7] = 4'h0;
    SS7[17][7] = 4'h0;
    SS7[18][7] = 4'h0;
    SS7[19][7] = 4'h0;
    SS7[20][7] = 4'h0;
    SS7[21][7] = 4'h0;
    SS7[22][7] = 4'h0;
    SS7[23][7] = 4'h0;
    SS7[24][7] = 4'hE;
    SS7[25][7] = 4'hD;
    SS7[26][7] = 4'hD;
    SS7[27][7] = 4'hC;
    SS7[28][7] = 4'hC;
    SS7[29][7] = 4'hC;
    SS7[30][7] = 4'h0;
    SS7[31][7] = 4'h0;
    SS7[32][7] = 4'h0;
    SS7[33][7] = 4'h0;
    SS7[34][7] = 4'h0;
    SS7[35][7] = 4'h0;
    SS7[36][7] = 4'h0;
    SS7[37][7] = 4'h0;
    SS7[38][7] = 4'h0;
    SS7[39][7] = 4'h0;
    SS7[40][7] = 4'h0;
    SS7[41][7] = 4'hD;
    SS7[42][7] = 4'hD;
    SS7[43][7] = 4'h0;
    SS7[44][7] = 4'h0;
    SS7[45][7] = 4'h0;
    SS7[46][7] = 4'h0;
    SS7[47][7] = 4'h0;
    SS7[0][8] = 4'h0;
    SS7[1][8] = 4'h0;
    SS7[2][8] = 4'hD;
    SS7[3][8] = 4'hD;
    SS7[4][8] = 4'hD;
    SS7[5][8] = 4'h0;
    SS7[6][8] = 4'h0;
    SS7[7][8] = 4'hD;
    SS7[8][8] = 4'h0;
    SS7[9][8] = 4'h0;
    SS7[10][8] = 4'h0;
    SS7[11][8] = 4'h0;
    SS7[12][8] = 4'h0;
    SS7[13][8] = 4'h0;
    SS7[14][8] = 4'h0;
    SS7[15][8] = 4'h0;
    SS7[16][8] = 4'h0;
    SS7[17][8] = 4'h0;
    SS7[18][8] = 4'h0;
    SS7[19][8] = 4'h0;
    SS7[20][8] = 4'h0;
    SS7[21][8] = 4'h0;
    SS7[22][8] = 4'h0;
    SS7[23][8] = 4'hE;
    SS7[24][8] = 4'hD;
    SS7[25][8] = 4'hD;
    SS7[26][8] = 4'hD;
    SS7[27][8] = 4'hC;
    SS7[28][8] = 4'hC;
    SS7[29][8] = 4'hC;
    SS7[30][8] = 4'h0;
    SS7[31][8] = 4'h0;
    SS7[32][8] = 4'h0;
    SS7[33][8] = 4'h0;
    SS7[34][8] = 4'h0;
    SS7[35][8] = 4'h0;
    SS7[36][8] = 4'h0;
    SS7[37][8] = 4'h0;
    SS7[38][8] = 4'hD;
    SS7[39][8] = 4'hD;
    SS7[40][8] = 4'hD;
    SS7[41][8] = 4'hD;
    SS7[42][8] = 4'hD;
    SS7[43][8] = 4'h0;
    SS7[44][8] = 4'h0;
    SS7[45][8] = 4'h0;
    SS7[46][8] = 4'h0;
    SS7[47][8] = 4'h0;
    SS7[0][9] = 4'h0;
    SS7[1][9] = 4'h0;
    SS7[2][9] = 4'hD;
    SS7[3][9] = 4'hD;
    SS7[4][9] = 4'hD;
    SS7[5][9] = 4'hD;
    SS7[6][9] = 4'hD;
    SS7[7][9] = 4'hD;
    SS7[8][9] = 4'h0;
    SS7[9][9] = 4'h0;
    SS7[10][9] = 4'h0;
    SS7[11][9] = 4'h0;
    SS7[12][9] = 4'h0;
    SS7[13][9] = 4'h0;
    SS7[14][9] = 4'h0;
    SS7[15][9] = 4'h0;
    SS7[16][9] = 4'h0;
    SS7[17][9] = 4'h0;
    SS7[18][9] = 4'h0;
    SS7[19][9] = 4'h0;
    SS7[20][9] = 4'h0;
    SS7[21][9] = 4'hE;
    SS7[22][9] = 4'hE;
    SS7[23][9] = 4'hE;
    SS7[24][9] = 4'hD;
    SS7[25][9] = 4'hD;
    SS7[26][9] = 4'hD;
    SS7[27][9] = 4'hD;
    SS7[28][9] = 4'hC;
    SS7[29][9] = 4'hC;
    SS7[30][9] = 4'hC;
    SS7[31][9] = 4'h0;
    SS7[32][9] = 4'h0;
    SS7[33][9] = 4'h0;
    SS7[34][9] = 4'h0;
    SS7[35][9] = 4'h0;
    SS7[36][9] = 4'hE;
    SS7[37][9] = 4'hD;
    SS7[38][9] = 4'hD;
    SS7[39][9] = 4'hD;
    SS7[40][9] = 4'hD;
    SS7[41][9] = 4'hD;
    SS7[42][9] = 4'hD;
    SS7[43][9] = 4'hD;
    SS7[44][9] = 4'h0;
    SS7[45][9] = 4'h0;
    SS7[46][9] = 4'h0;
    SS7[47][9] = 4'h0;
    SS7[0][10] = 4'h0;
    SS7[1][10] = 4'h0;
    SS7[2][10] = 4'hC;
    SS7[3][10] = 4'hC;
    SS7[4][10] = 4'hC;
    SS7[5][10] = 4'hC;
    SS7[6][10] = 4'hD;
    SS7[7][10] = 4'hD;
    SS7[8][10] = 4'hD;
    SS7[9][10] = 4'h0;
    SS7[10][10] = 4'hE;
    SS7[11][10] = 4'hE;
    SS7[12][10] = 4'h0;
    SS7[13][10] = 4'h0;
    SS7[14][10] = 4'h0;
    SS7[15][10] = 4'h0;
    SS7[16][10] = 4'h0;
    SS7[17][10] = 4'h0;
    SS7[18][10] = 4'h0;
    SS7[19][10] = 4'h0;
    SS7[20][10] = 4'h0;
    SS7[21][10] = 4'h0;
    SS7[22][10] = 4'hE;
    SS7[23][10] = 4'hE;
    SS7[24][10] = 4'hE;
    SS7[25][10] = 4'hD;
    SS7[26][10] = 4'hC;
    SS7[27][10] = 4'hC;
    SS7[28][10] = 4'hC;
    SS7[29][10] = 4'hC;
    SS7[30][10] = 4'hC;
    SS7[31][10] = 4'h0;
    SS7[32][10] = 4'h0;
    SS7[33][10] = 4'hE;
    SS7[34][10] = 4'hE;
    SS7[35][10] = 4'hE;
    SS7[36][10] = 4'hE;
    SS7[37][10] = 4'hE;
    SS7[38][10] = 4'hD;
    SS7[39][10] = 4'hD;
    SS7[40][10] = 4'hD;
    SS7[41][10] = 4'h0;
    SS7[42][10] = 4'h0;
    SS7[43][10] = 4'h0;
    SS7[44][10] = 4'h0;
    SS7[45][10] = 4'h0;
    SS7[46][10] = 4'h0;
    SS7[47][10] = 4'h0;
    SS7[0][11] = 4'h0;
    SS7[1][11] = 4'h0;
    SS7[2][11] = 4'h0;
    SS7[3][11] = 4'hC;
    SS7[4][11] = 4'hC;
    SS7[5][11] = 4'hC;
    SS7[6][11] = 4'hD;
    SS7[7][11] = 4'hD;
    SS7[8][11] = 4'hC;
    SS7[9][11] = 4'hE;
    SS7[10][11] = 4'hE;
    SS7[11][11] = 4'hE;
    SS7[12][11] = 4'h0;
    SS7[13][11] = 4'h0;
    SS7[14][11] = 4'h0;
    SS7[15][11] = 4'hE;
    SS7[16][11] = 4'h0;
    SS7[17][11] = 4'h0;
    SS7[18][11] = 4'h0;
    SS7[19][11] = 4'h0;
    SS7[20][11] = 4'h0;
    SS7[21][11] = 4'h0;
    SS7[22][11] = 4'hE;
    SS7[23][11] = 4'hD;
    SS7[24][11] = 4'hD;
    SS7[25][11] = 4'hC;
    SS7[26][11] = 4'hC;
    SS7[27][11] = 4'hC;
    SS7[28][11] = 4'hC;
    SS7[29][11] = 4'hC;
    SS7[30][11] = 4'hC;
    SS7[31][11] = 4'hC;
    SS7[32][11] = 4'hE;
    SS7[33][11] = 4'hE;
    SS7[34][11] = 4'hE;
    SS7[35][11] = 4'hE;
    SS7[36][11] = 4'hE;
    SS7[37][11] = 4'hE;
    SS7[38][11] = 4'hD;
    SS7[39][11] = 4'hD;
    SS7[40][11] = 4'hD;
    SS7[41][11] = 4'h0;
    SS7[42][11] = 4'h0;
    SS7[43][11] = 4'h0;
    SS7[44][11] = 4'h0;
    SS7[45][11] = 4'h0;
    SS7[46][11] = 4'h0;
    SS7[47][11] = 4'h0;
    SS7[0][12] = 4'h0;
    SS7[1][12] = 4'h0;
    SS7[2][12] = 4'h0;
    SS7[3][12] = 4'hC;
    SS7[4][12] = 4'hC;
    SS7[5][12] = 4'hC;
    SS7[6][12] = 4'hC;
    SS7[7][12] = 4'hC;
    SS7[8][12] = 4'hC;
    SS7[9][12] = 4'hC;
    SS7[10][12] = 4'hE;
    SS7[11][12] = 4'hE;
    SS7[12][12] = 4'hE;
    SS7[13][12] = 4'hE;
    SS7[14][12] = 4'hE;
    SS7[15][12] = 4'hE;
    SS7[16][12] = 4'h0;
    SS7[17][12] = 4'h0;
    SS7[18][12] = 4'h0;
    SS7[19][12] = 4'h0;
    SS7[20][12] = 4'h0;
    SS7[21][12] = 4'hE;
    SS7[22][12] = 4'hD;
    SS7[23][12] = 4'hD;
    SS7[24][12] = 4'hD;
    SS7[25][12] = 4'hD;
    SS7[26][12] = 4'hC;
    SS7[27][12] = 4'hC;
    SS7[28][12] = 4'hC;
    SS7[29][12] = 4'hC;
    SS7[30][12] = 4'hC;
    SS7[31][12] = 4'hC;
    SS7[32][12] = 4'hE;
    SS7[33][12] = 4'hE;
    SS7[34][12] = 4'hE;
    SS7[35][12] = 4'hE;
    SS7[36][12] = 4'hD;
    SS7[37][12] = 4'hD;
    SS7[38][12] = 4'hD;
    SS7[39][12] = 4'hD;
    SS7[40][12] = 4'hD;
    SS7[41][12] = 4'hD;
    SS7[42][12] = 4'h0;
    SS7[43][12] = 4'h0;
    SS7[44][12] = 4'h0;
    SS7[45][12] = 4'h0;
    SS7[46][12] = 4'h0;
    SS7[47][12] = 4'h0;
    SS7[0][13] = 4'h0;
    SS7[1][13] = 4'h0;
    SS7[2][13] = 4'h0;
    SS7[3][13] = 4'h0;
    SS7[4][13] = 4'hC;
    SS7[5][13] = 4'hC;
    SS7[6][13] = 4'hC;
    SS7[7][13] = 4'hC;
    SS7[8][13] = 4'hC;
    SS7[9][13] = 4'hC;
    SS7[10][13] = 4'hE;
    SS7[11][13] = 4'hD;
    SS7[12][13] = 4'hD;
    SS7[13][13] = 4'hE;
    SS7[14][13] = 4'hE;
    SS7[15][13] = 4'hE;
    SS7[16][13] = 4'h0;
    SS7[17][13] = 4'h0;
    SS7[18][13] = 4'hE;
    SS7[19][13] = 4'hE;
    SS7[20][13] = 4'hE;
    SS7[21][13] = 4'hE;
    SS7[22][13] = 4'hE;
    SS7[23][13] = 4'hD;
    SS7[24][13] = 4'hD;
    SS7[25][13] = 4'hD;
    SS7[26][13] = 4'hC;
    SS7[27][13] = 4'hC;
    SS7[28][13] = 4'hC;
    SS7[29][13] = 4'hC;
    SS7[30][13] = 4'hC;
    SS7[31][13] = 4'hC;
    SS7[32][13] = 4'hE;
    SS7[33][13] = 4'hE;
    SS7[34][13] = 4'hE;
    SS7[35][13] = 4'hE;
    SS7[36][13] = 4'hD;
    SS7[37][13] = 4'hD;
    SS7[38][13] = 4'hD;
    SS7[39][13] = 4'hD;
    SS7[40][13] = 4'hD;
    SS7[41][13] = 4'hD;
    SS7[42][13] = 4'h0;
    SS7[43][13] = 4'h0;
    SS7[44][13] = 4'h0;
    SS7[45][13] = 4'h0;
    SS7[46][13] = 4'h0;
    SS7[47][13] = 4'h0;
    SS7[0][14] = 4'h0;
    SS7[1][14] = 4'h0;
    SS7[2][14] = 4'h0;
    SS7[3][14] = 4'h0;
    SS7[4][14] = 4'hC;
    SS7[5][14] = 4'hC;
    SS7[6][14] = 4'hC;
    SS7[7][14] = 4'hC;
    SS7[8][14] = 4'hC;
    SS7[9][14] = 4'hC;
    SS7[10][14] = 4'hD;
    SS7[11][14] = 4'hD;
    SS7[12][14] = 4'hD;
    SS7[13][14] = 4'hD;
    SS7[14][14] = 4'hE;
    SS7[15][14] = 4'hE;
    SS7[16][14] = 4'hD;
    SS7[17][14] = 4'hE;
    SS7[18][14] = 4'hE;
    SS7[19][14] = 4'hE;
    SS7[20][14] = 4'hE;
    SS7[21][14] = 4'hE;
    SS7[22][14] = 4'hE;
    SS7[23][14] = 4'hD;
    SS7[24][14] = 4'hC;
    SS7[25][14] = 4'hC;
    SS7[26][14] = 4'hC;
    SS7[27][14] = 4'hC;
    SS7[28][14] = 4'hC;
    SS7[29][14] = 4'hC;
    SS7[30][14] = 4'hC;
    SS7[31][14] = 4'hE;
    SS7[32][14] = 4'hE;
    SS7[33][14] = 4'hE;
    SS7[34][14] = 4'hE;
    SS7[35][14] = 4'hE;
    SS7[36][14] = 4'hD;
    SS7[37][14] = 4'hD;
    SS7[38][14] = 4'hD;
    SS7[39][14] = 4'h0;
    SS7[40][14] = 4'h0;
    SS7[41][14] = 4'h0;
    SS7[42][14] = 4'h0;
    SS7[43][14] = 4'h0;
    SS7[44][14] = 4'h0;
    SS7[45][14] = 4'h0;
    SS7[46][14] = 4'h0;
    SS7[47][14] = 4'h0;
    SS7[0][15] = 4'h0;
    SS7[1][15] = 4'h0;
    SS7[2][15] = 4'h0;
    SS7[3][15] = 4'h0;
    SS7[4][15] = 4'hC;
    SS7[5][15] = 4'hC;
    SS7[6][15] = 4'h0;
    SS7[7][15] = 4'h0;
    SS7[8][15] = 4'hC;
    SS7[9][15] = 4'hC;
    SS7[10][15] = 4'hC;
    SS7[11][15] = 4'hD;
    SS7[12][15] = 4'hD;
    SS7[13][15] = 4'hD;
    SS7[14][15] = 4'hD;
    SS7[15][15] = 4'hD;
    SS7[16][15] = 4'hD;
    SS7[17][15] = 4'hE;
    SS7[18][15] = 4'hE;
    SS7[19][15] = 4'hE;
    SS7[20][15] = 4'hE;
    SS7[21][15] = 4'hE;
    SS7[22][15] = 4'hE;
    SS7[23][15] = 4'hE;
    SS7[24][15] = 4'hC;
    SS7[25][15] = 4'hC;
    SS7[26][15] = 4'hC;
    SS7[27][15] = 4'hC;
    SS7[28][15] = 4'hC;
    SS7[29][15] = 4'hC;
    SS7[30][15] = 4'hE;
    SS7[31][15] = 4'hE;
    SS7[32][15] = 4'hE;
    SS7[33][15] = 4'hE;
    SS7[34][15] = 4'hE;
    SS7[35][15] = 4'hE;
    SS7[36][15] = 4'hE;
    SS7[37][15] = 4'h3;
    SS7[38][15] = 4'h3;
    SS7[39][15] = 4'h3;
    SS7[40][15] = 4'h0;
    SS7[41][15] = 4'h0;
    SS7[42][15] = 4'h0;
    SS7[43][15] = 4'h0;
    SS7[44][15] = 4'h0;
    SS7[45][15] = 4'h0;
    SS7[46][15] = 4'h0;
    SS7[47][15] = 4'h0;
    SS7[0][16] = 4'h0;
    SS7[1][16] = 4'h0;
    SS7[2][16] = 4'h0;
    SS7[3][16] = 4'h0;
    SS7[4][16] = 4'h0;
    SS7[5][16] = 4'h0;
    SS7[6][16] = 4'h0;
    SS7[7][16] = 4'h0;
    SS7[8][16] = 4'hC;
    SS7[9][16] = 4'hC;
    SS7[10][16] = 4'hC;
    SS7[11][16] = 4'hC;
    SS7[12][16] = 4'hC;
    SS7[13][16] = 4'hC;
    SS7[14][16] = 4'hD;
    SS7[15][16] = 4'hD;
    SS7[16][16] = 4'hD;
    SS7[17][16] = 4'hD;
    SS7[18][16] = 4'hE;
    SS7[19][16] = 4'hE;
    SS7[20][16] = 4'hE;
    SS7[21][16] = 4'hE;
    SS7[22][16] = 4'hE;
    SS7[23][16] = 4'hE;
    SS7[24][16] = 4'hC;
    SS7[25][16] = 4'hC;
    SS7[26][16] = 4'hC;
    SS7[27][16] = 4'hC;
    SS7[28][16] = 4'hC;
    SS7[29][16] = 4'hC;
    SS7[30][16] = 4'hC;
    SS7[31][16] = 4'hE;
    SS7[32][16] = 4'hE;
    SS7[33][16] = 4'hE;
    SS7[34][16] = 4'hD;
    SS7[35][16] = 4'hD;
    SS7[36][16] = 4'hD;
    SS7[37][16] = 4'h3;
    SS7[38][16] = 4'h3;
    SS7[39][16] = 4'h3;
    SS7[40][16] = 4'h0;
    SS7[41][16] = 4'h0;
    SS7[42][16] = 4'h0;
    SS7[43][16] = 4'h0;
    SS7[44][16] = 4'h0;
    SS7[45][16] = 4'h0;
    SS7[46][16] = 4'h0;
    SS7[47][16] = 4'h0;
    SS7[0][17] = 4'h0;
    SS7[1][17] = 4'h0;
    SS7[2][17] = 4'h0;
    SS7[3][17] = 4'h0;
    SS7[4][17] = 4'h0;
    SS7[5][17] = 4'h0;
    SS7[6][17] = 4'h0;
    SS7[7][17] = 4'h0;
    SS7[8][17] = 4'hC;
    SS7[9][17] = 4'hC;
    SS7[10][17] = 4'hC;
    SS7[11][17] = 4'hC;
    SS7[12][17] = 4'hC;
    SS7[13][17] = 4'hC;
    SS7[14][17] = 4'hC;
    SS7[15][17] = 4'hD;
    SS7[16][17] = 4'hC;
    SS7[17][17] = 4'hC;
    SS7[18][17] = 4'hE;
    SS7[19][17] = 4'hE;
    SS7[20][17] = 4'hE;
    SS7[21][17] = 4'hE;
    SS7[22][17] = 4'hE;
    SS7[23][17] = 4'hE;
    SS7[24][17] = 4'hD;
    SS7[25][17] = 4'hC;
    SS7[26][17] = 4'hC;
    SS7[27][17] = 4'hC;
    SS7[28][17] = 4'hC;
    SS7[29][17] = 4'hC;
    SS7[30][17] = 4'hC;
    SS7[31][17] = 4'hE;
    SS7[32][17] = 4'hD;
    SS7[33][17] = 4'hD;
    SS7[34][17] = 4'hD;
    SS7[35][17] = 4'hD;
    SS7[36][17] = 4'hD;
    SS7[37][17] = 4'h3;
    SS7[38][17] = 4'h3;
    SS7[39][17] = 4'h3;
    SS7[40][17] = 4'h0;
    SS7[41][17] = 4'h0;
    SS7[42][17] = 4'h0;
    SS7[43][17] = 4'h0;
    SS7[44][17] = 4'h0;
    SS7[45][17] = 4'h0;
    SS7[46][17] = 4'h0;
    SS7[47][17] = 4'h0;
    SS7[0][18] = 4'h0;
    SS7[1][18] = 4'h0;
    SS7[2][18] = 4'h0;
    SS7[3][18] = 4'h0;
    SS7[4][18] = 4'h0;
    SS7[5][18] = 4'h0;
    SS7[6][18] = 4'h0;
    SS7[7][18] = 4'h0;
    SS7[8][18] = 4'h0;
    SS7[9][18] = 4'hC;
    SS7[10][18] = 4'hC;
    SS7[11][18] = 4'hC;
    SS7[12][18] = 4'hC;
    SS7[13][18] = 4'hC;
    SS7[14][18] = 4'hC;
    SS7[15][18] = 4'hC;
    SS7[16][18] = 4'hC;
    SS7[17][18] = 4'hC;
    SS7[18][18] = 4'hC;
    SS7[19][18] = 4'hE;
    SS7[20][18] = 4'hE;
    SS7[21][18] = 4'hE;
    SS7[22][18] = 4'hD;
    SS7[23][18] = 4'hD;
    SS7[24][18] = 4'hD;
    SS7[25][18] = 4'hC;
    SS7[26][18] = 4'hC;
    SS7[27][18] = 4'hC;
    SS7[28][18] = 4'hC;
    SS7[29][18] = 4'hC;
    SS7[30][18] = 4'hE;
    SS7[31][18] = 4'hD;
    SS7[32][18] = 4'hD;
    SS7[33][18] = 4'hD;
    SS7[34][18] = 4'hD;
    SS7[35][18] = 4'hD;
    SS7[36][18] = 4'hD;
    SS7[37][18] = 4'h0;
    SS7[38][18] = 4'h0;
    SS7[39][18] = 4'h0;
    SS7[40][18] = 4'h0;
    SS7[41][18] = 4'h0;
    SS7[42][18] = 4'h0;
    SS7[43][18] = 4'h0;
    SS7[44][18] = 4'h0;
    SS7[45][18] = 4'h0;
    SS7[46][18] = 4'h0;
    SS7[47][18] = 4'h0;
    SS7[0][19] = 4'h0;
    SS7[1][19] = 4'h0;
    SS7[2][19] = 4'h0;
    SS7[3][19] = 4'h0;
    SS7[4][19] = 4'h0;
    SS7[5][19] = 4'h0;
    SS7[6][19] = 4'h0;
    SS7[7][19] = 4'h0;
    SS7[8][19] = 4'h0;
    SS7[9][19] = 4'hC;
    SS7[10][19] = 4'hC;
    SS7[11][19] = 4'hC;
    SS7[12][19] = 4'hC;
    SS7[13][19] = 4'hC;
    SS7[14][19] = 4'hC;
    SS7[15][19] = 4'hC;
    SS7[16][19] = 4'hC;
    SS7[17][19] = 4'hC;
    SS7[18][19] = 4'hC;
    SS7[19][19] = 4'hD;
    SS7[20][19] = 4'hD;
    SS7[21][19] = 4'hD;
    SS7[22][19] = 4'hD;
    SS7[23][19] = 4'hD;
    SS7[24][19] = 4'hD;
    SS7[25][19] = 4'hC;
    SS7[26][19] = 4'hC;
    SS7[27][19] = 4'hC;
    SS7[28][19] = 4'hC;
    SS7[29][19] = 4'hE;
    SS7[30][19] = 4'hE;
    SS7[31][19] = 4'hE;
    SS7[32][19] = 4'hD;
    SS7[33][19] = 4'hD;
    SS7[34][19] = 4'hD;
    SS7[35][19] = 4'h0;
    SS7[36][19] = 4'h0;
    SS7[37][19] = 4'h0;
    SS7[38][19] = 4'h0;
    SS7[39][19] = 4'h0;
    SS7[40][19] = 4'h0;
    SS7[41][19] = 4'h0;
    SS7[42][19] = 4'h0;
    SS7[43][19] = 4'h0;
    SS7[44][19] = 4'h0;
    SS7[45][19] = 4'h0;
    SS7[46][19] = 4'h0;
    SS7[47][19] = 4'h0;
    SS7[0][20] = 4'h0;
    SS7[1][20] = 4'h0;
    SS7[2][20] = 4'h0;
    SS7[3][20] = 4'h0;
    SS7[4][20] = 4'h0;
    SS7[5][20] = 4'h0;
    SS7[6][20] = 4'h0;
    SS7[7][20] = 4'h0;
    SS7[8][20] = 4'h0;
    SS7[9][20] = 4'hE;
    SS7[10][20] = 4'hC;
    SS7[11][20] = 4'hC;
    SS7[12][20] = 4'hC;
    SS7[13][20] = 4'hC;
    SS7[14][20] = 4'hC;
    SS7[15][20] = 4'hC;
    SS7[16][20] = 4'hC;
    SS7[17][20] = 4'hC;
    SS7[18][20] = 4'hC;
    SS7[19][20] = 4'hD;
    SS7[20][20] = 4'hD;
    SS7[21][20] = 4'hD;
    SS7[22][20] = 4'hD;
    SS7[23][20] = 4'hD;
    SS7[24][20] = 4'hD;
    SS7[25][20] = 4'hC;
    SS7[26][20] = 4'hC;
    SS7[27][20] = 4'hC;
    SS7[28][20] = 4'hC;
    SS7[29][20] = 4'hE;
    SS7[30][20] = 4'hE;
    SS7[31][20] = 4'hE;
    SS7[32][20] = 4'hD;
    SS7[33][20] = 4'hD;
    SS7[34][20] = 4'hD;
    SS7[35][20] = 4'h0;
    SS7[36][20] = 4'h0;
    SS7[37][20] = 4'h0;
    SS7[38][20] = 4'h0;
    SS7[39][20] = 4'h0;
    SS7[40][20] = 4'h0;
    SS7[41][20] = 4'h0;
    SS7[42][20] = 4'h0;
    SS7[43][20] = 4'h0;
    SS7[44][20] = 4'h0;
    SS7[45][20] = 4'h0;
    SS7[46][20] = 4'h0;
    SS7[47][20] = 4'h0;
    SS7[0][21] = 4'h0;
    SS7[1][21] = 4'h0;
    SS7[2][21] = 4'h0;
    SS7[3][21] = 4'h0;
    SS7[4][21] = 4'h0;
    SS7[5][21] = 4'h0;
    SS7[6][21] = 4'h0;
    SS7[7][21] = 4'hE;
    SS7[8][21] = 4'hE;
    SS7[9][21] = 4'hE;
    SS7[10][21] = 4'hC;
    SS7[11][21] = 4'hC;
    SS7[12][21] = 4'hC;
    SS7[13][21] = 4'hC;
    SS7[14][21] = 4'hC;
    SS7[15][21] = 4'hC;
    SS7[16][21] = 4'hC;
    SS7[17][21] = 4'hC;
    SS7[18][21] = 4'hC;
    SS7[19][21] = 4'hC;
    SS7[20][21] = 4'hD;
    SS7[21][21] = 4'hD;
    SS7[22][21] = 4'hC;
    SS7[23][21] = 4'hC;
    SS7[24][21] = 4'hC;
    SS7[25][21] = 4'hC;
    SS7[26][21] = 4'hC;
    SS7[27][21] = 4'hC;
    SS7[28][21] = 4'hC;
    SS7[29][21] = 4'hE;
    SS7[30][21] = 4'hD;
    SS7[31][21] = 4'hD;
    SS7[32][21] = 4'hD;
    SS7[33][21] = 4'hD;
    SS7[34][21] = 4'hD;
    SS7[35][21] = 4'hD;
    SS7[36][21] = 4'h0;
    SS7[37][21] = 4'h0;
    SS7[38][21] = 4'h0;
    SS7[39][21] = 4'h0;
    SS7[40][21] = 4'h0;
    SS7[41][21] = 4'h0;
    SS7[42][21] = 4'h0;
    SS7[43][21] = 4'h0;
    SS7[44][21] = 4'h0;
    SS7[45][21] = 4'h0;
    SS7[46][21] = 4'h0;
    SS7[47][21] = 4'h0;
    SS7[0][22] = 4'h0;
    SS7[1][22] = 4'h0;
    SS7[2][22] = 4'h0;
    SS7[3][22] = 4'h0;
    SS7[4][22] = 4'hE;
    SS7[5][22] = 4'hE;
    SS7[6][22] = 4'hE;
    SS7[7][22] = 4'hE;
    SS7[8][22] = 4'hE;
    SS7[9][22] = 4'hE;
    SS7[10][22] = 4'hE;
    SS7[11][22] = 4'hC;
    SS7[12][22] = 4'hE;
    SS7[13][22] = 4'hE;
    SS7[14][22] = 4'hC;
    SS7[15][22] = 4'hC;
    SS7[16][22] = 4'hC;
    SS7[17][22] = 4'hC;
    SS7[18][22] = 4'hC;
    SS7[19][22] = 4'hC;
    SS7[20][22] = 4'hC;
    SS7[21][22] = 4'hC;
    SS7[22][22] = 4'hC;
    SS7[23][22] = 4'hC;
    SS7[24][22] = 4'hC;
    SS7[25][22] = 4'hC;
    SS7[26][22] = 4'hC;
    SS7[27][22] = 4'hC;
    SS7[28][22] = 4'hC;
    SS7[29][22] = 4'hC;
    SS7[30][22] = 4'hD;
    SS7[31][22] = 4'hD;
    SS7[32][22] = 4'hD;
    SS7[33][22] = 4'hD;
    SS7[34][22] = 4'hD;
    SS7[35][22] = 4'h3;
    SS7[36][22] = 4'h0;
    SS7[37][22] = 4'h0;
    SS7[38][22] = 4'h0;
    SS7[39][22] = 4'h0;
    SS7[40][22] = 4'h0;
    SS7[41][22] = 4'h0;
    SS7[42][22] = 4'h0;
    SS7[43][22] = 4'h0;
    SS7[44][22] = 4'h0;
    SS7[45][22] = 4'h0;
    SS7[46][22] = 4'h0;
    SS7[47][22] = 4'h0;
    SS7[0][23] = 4'h0;
    SS7[1][23] = 4'h0;
    SS7[2][23] = 4'hD;
    SS7[3][23] = 4'hD;
    SS7[4][23] = 4'hD;
    SS7[5][23] = 4'hE;
    SS7[6][23] = 4'hE;
    SS7[7][23] = 4'hE;
    SS7[8][23] = 4'hE;
    SS7[9][23] = 4'hE;
    SS7[10][23] = 4'hE;
    SS7[11][23] = 4'hE;
    SS7[12][23] = 4'hE;
    SS7[13][23] = 4'hE;
    SS7[14][23] = 4'hC;
    SS7[15][23] = 4'hC;
    SS7[16][23] = 4'hC;
    SS7[17][23] = 4'hC;
    SS7[18][23] = 4'hC;
    SS7[19][23] = 4'hC;
    SS7[20][23] = 4'hC;
    SS7[21][23] = 4'hC;
    SS7[22][23] = 4'hC;
    SS7[23][23] = 4'hC;
    SS7[24][23] = 4'hC;
    SS7[25][23] = 4'hD;
    SS7[26][23] = 4'hD;
    SS7[27][23] = 4'hC;
    SS7[28][23] = 4'hC;
    SS7[29][23] = 4'hC;
    SS7[30][23] = 4'hD;
    SS7[31][23] = 4'hD;
    SS7[32][23] = 4'hD;
    SS7[33][23] = 4'h3;
    SS7[34][23] = 4'h3;
    SS7[35][23] = 4'h3;
    SS7[36][23] = 4'h3;
    SS7[37][23] = 4'h0;
    SS7[38][23] = 4'h0;
    SS7[39][23] = 4'h0;
    SS7[40][23] = 4'h0;
    SS7[41][23] = 4'h0;
    SS7[42][23] = 4'h0;
    SS7[43][23] = 4'h0;
    SS7[44][23] = 4'h0;
    SS7[45][23] = 4'h0;
    SS7[46][23] = 4'h0;
    SS7[47][23] = 4'h0;
    SS7[0][24] = 4'hD;
    SS7[1][24] = 4'hD;
    SS7[2][24] = 4'hD;
    SS7[3][24] = 4'hD;
    SS7[4][24] = 4'hD;
    SS7[5][24] = 4'hE;
    SS7[6][24] = 4'hE;
    SS7[7][24] = 4'hD;
    SS7[8][24] = 4'hE;
    SS7[9][24] = 4'hE;
    SS7[10][24] = 4'hE;
    SS7[11][24] = 4'hE;
    SS7[12][24] = 4'hE;
    SS7[13][24] = 4'hE;
    SS7[14][24] = 4'hE;
    SS7[15][24] = 4'hE;
    SS7[16][24] = 4'hE;
    SS7[17][24] = 4'hE;
    SS7[18][24] = 4'hC;
    SS7[19][24] = 4'hC;
    SS7[20][24] = 4'hC;
    SS7[21][24] = 4'hC;
    SS7[22][24] = 4'hC;
    SS7[23][24] = 4'hD;
    SS7[24][24] = 4'hD;
    SS7[25][24] = 4'hD;
    SS7[26][24] = 4'hD;
    SS7[27][24] = 4'hC;
    SS7[28][24] = 4'hC;
    SS7[29][24] = 4'hC;
    SS7[30][24] = 4'hC;
    SS7[31][24] = 4'hD;
    SS7[32][24] = 4'hD;
    SS7[33][24] = 4'hD;
    SS7[34][24] = 4'h3;
    SS7[35][24] = 4'h3;
    SS7[36][24] = 4'h3;
    SS7[37][24] = 4'h0;
    SS7[38][24] = 4'h0;
    SS7[39][24] = 4'h0;
    SS7[40][24] = 4'h0;
    SS7[41][24] = 4'h0;
    SS7[42][24] = 4'h0;
    SS7[43][24] = 4'h0;
    SS7[44][24] = 4'h0;
    SS7[45][24] = 4'h0;
    SS7[46][24] = 4'h0;
    SS7[47][24] = 4'h0;
    SS7[0][25] = 4'hD;
    SS7[1][25] = 4'hD;
    SS7[2][25] = 4'hD;
    SS7[3][25] = 4'hD;
    SS7[4][25] = 4'hD;
    SS7[5][25] = 4'hD;
    SS7[6][25] = 4'hD;
    SS7[7][25] = 4'hD;
    SS7[8][25] = 4'hD;
    SS7[9][25] = 4'hE;
    SS7[10][25] = 4'hE;
    SS7[11][25] = 4'hE;
    SS7[12][25] = 4'hE;
    SS7[13][25] = 4'hD;
    SS7[14][25] = 4'hD;
    SS7[15][25] = 4'hE;
    SS7[16][25] = 4'hE;
    SS7[17][25] = 4'hE;
    SS7[18][25] = 4'hC;
    SS7[19][25] = 4'hC;
    SS7[20][25] = 4'hC;
    SS7[21][25] = 4'hD;
    SS7[22][25] = 4'hD;
    SS7[23][25] = 4'hD;
    SS7[24][25] = 4'hD;
    SS7[25][25] = 4'hD;
    SS7[26][25] = 4'hD;
    SS7[27][25] = 4'hD;
    SS7[28][25] = 4'hD;
    SS7[29][25] = 4'hD;
    SS7[30][25] = 4'hD;
    SS7[31][25] = 4'hD;
    SS7[32][25] = 4'hD;
    SS7[33][25] = 4'hD;
    SS7[34][25] = 4'h3;
    SS7[35][25] = 4'h3;
    SS7[36][25] = 4'h0;
    SS7[37][25] = 4'h0;
    SS7[38][25] = 4'h0;
    SS7[39][25] = 4'h0;
    SS7[40][25] = 4'h0;
    SS7[41][25] = 4'h0;
    SS7[42][25] = 4'h0;
    SS7[43][25] = 4'h0;
    SS7[44][25] = 4'h0;
    SS7[45][25] = 4'h0;
    SS7[46][25] = 4'h0;
    SS7[47][25] = 4'h0;
    SS7[0][26] = 4'hD;
    SS7[1][26] = 4'hD;
    SS7[2][26] = 4'hE;
    SS7[3][26] = 4'hD;
    SS7[4][26] = 4'hD;
    SS7[5][26] = 4'hD;
    SS7[6][26] = 4'hD;
    SS7[7][26] = 4'hD;
    SS7[8][26] = 4'hD;
    SS7[9][26] = 4'hE;
    SS7[10][26] = 4'hD;
    SS7[11][26] = 4'hD;
    SS7[12][26] = 4'hD;
    SS7[13][26] = 4'hD;
    SS7[14][26] = 4'hD;
    SS7[15][26] = 4'hE;
    SS7[16][26] = 4'hE;
    SS7[17][26] = 4'hE;
    SS7[18][26] = 4'hD;
    SS7[19][26] = 4'hC;
    SS7[20][26] = 4'hC;
    SS7[21][26] = 4'hC;
    SS7[22][26] = 4'hD;
    SS7[23][26] = 4'hD;
    SS7[24][26] = 4'hD;
    SS7[25][26] = 4'hD;
    SS7[26][26] = 4'hA;
    SS7[27][26] = 4'hA;
    SS7[28][26] = 4'hD;
    SS7[29][26] = 4'hD;
    SS7[30][26] = 4'hD;
    SS7[31][26] = 4'hD;
    SS7[32][26] = 4'hD;
    SS7[33][26] = 4'hF;
    SS7[34][26] = 4'h0;
    SS7[35][26] = 4'h0;
    SS7[36][26] = 4'h0;
    SS7[37][26] = 4'h0;
    SS7[38][26] = 4'h0;
    SS7[39][26] = 4'h0;
    SS7[40][26] = 4'h0;
    SS7[41][26] = 4'h0;
    SS7[42][26] = 4'h0;
    SS7[43][26] = 4'h0;
    SS7[44][26] = 4'h0;
    SS7[45][26] = 4'h0;
    SS7[46][26] = 4'h0;
    SS7[47][26] = 4'h0;
    SS7[0][27] = 4'h0;
    SS7[1][27] = 4'h0;
    SS7[2][27] = 4'h0;
    SS7[3][27] = 4'hD;
    SS7[4][27] = 4'hD;
    SS7[5][27] = 4'hD;
    SS7[6][27] = 4'hD;
    SS7[7][27] = 4'hD;
    SS7[8][27] = 4'h3;
    SS7[9][27] = 4'hD;
    SS7[10][27] = 4'hD;
    SS7[11][27] = 4'hD;
    SS7[12][27] = 4'hD;
    SS7[13][27] = 4'hD;
    SS7[14][27] = 4'hD;
    SS7[15][27] = 4'hD;
    SS7[16][27] = 4'hD;
    SS7[17][27] = 4'hD;
    SS7[18][27] = 4'hD;
    SS7[19][27] = 4'hC;
    SS7[20][27] = 4'hC;
    SS7[21][27] = 4'hC;
    SS7[22][27] = 4'hD;
    SS7[23][27] = 4'hA;
    SS7[24][27] = 4'hA;
    SS7[25][27] = 4'hA;
    SS7[26][27] = 4'hA;
    SS7[27][27] = 4'hA;
    SS7[28][27] = 4'hA;
    SS7[29][27] = 4'hD;
    SS7[30][27] = 4'hD;
    SS7[31][27] = 4'hC;
    SS7[32][27] = 4'h0;
    SS7[33][27] = 4'h0;
    SS7[34][27] = 4'h0;
    SS7[35][27] = 4'h0;
    SS7[36][27] = 4'h0;
    SS7[37][27] = 4'h0;
    SS7[38][27] = 4'h0;
    SS7[39][27] = 4'h0;
    SS7[40][27] = 4'h0;
    SS7[41][27] = 4'h0;
    SS7[42][27] = 4'h0;
    SS7[43][27] = 4'h0;
    SS7[44][27] = 4'h0;
    SS7[45][27] = 4'h0;
    SS7[46][27] = 4'h0;
    SS7[47][27] = 4'h0;
    SS7[0][28] = 4'h0;
    SS7[1][28] = 4'h0;
    SS7[2][28] = 4'h0;
    SS7[3][28] = 4'hD;
    SS7[4][28] = 4'hD;
    SS7[5][28] = 4'h0;
    SS7[6][28] = 4'h0;
    SS7[7][28] = 4'h3;
    SS7[8][28] = 4'h3;
    SS7[9][28] = 4'h3;
    SS7[10][28] = 4'hD;
    SS7[11][28] = 4'hD;
    SS7[12][28] = 4'hD;
    SS7[13][28] = 4'hD;
    SS7[14][28] = 4'hD;
    SS7[15][28] = 4'hD;
    SS7[16][28] = 4'hD;
    SS7[17][28] = 4'hD;
    SS7[18][28] = 4'hD;
    SS7[19][28] = 4'hC;
    SS7[20][28] = 4'hC;
    SS7[21][28] = 4'hD;
    SS7[22][28] = 4'hD;
    SS7[23][28] = 4'hA;
    SS7[24][28] = 4'hA;
    SS7[25][28] = 4'hA;
    SS7[26][28] = 4'hA;
    SS7[27][28] = 4'hA;
    SS7[28][28] = 4'hA;
    SS7[29][28] = 4'hC;
    SS7[30][28] = 4'hC;
    SS7[31][28] = 4'hC;
    SS7[32][28] = 4'h0;
    SS7[33][28] = 4'h0;
    SS7[34][28] = 4'h0;
    SS7[35][28] = 4'h0;
    SS7[36][28] = 4'h0;
    SS7[37][28] = 4'h0;
    SS7[38][28] = 4'h0;
    SS7[39][28] = 4'h0;
    SS7[40][28] = 4'h0;
    SS7[41][28] = 4'h0;
    SS7[42][28] = 4'h0;
    SS7[43][28] = 4'h0;
    SS7[44][28] = 4'h0;
    SS7[45][28] = 4'h0;
    SS7[46][28] = 4'h0;
    SS7[47][28] = 4'h0;
    SS7[0][29] = 4'h0;
    SS7[1][29] = 4'h0;
    SS7[2][29] = 4'h0;
    SS7[3][29] = 4'h0;
    SS7[4][29] = 4'h0;
    SS7[5][29] = 4'h0;
    SS7[6][29] = 4'h0;
    SS7[7][29] = 4'h3;
    SS7[8][29] = 4'h3;
    SS7[9][29] = 4'h3;
    SS7[10][29] = 4'hD;
    SS7[11][29] = 4'h0;
    SS7[12][29] = 4'h0;
    SS7[13][29] = 4'hD;
    SS7[14][29] = 4'hD;
    SS7[15][29] = 4'hD;
    SS7[16][29] = 4'hD;
    SS7[17][29] = 4'hD;
    SS7[18][29] = 4'hD;
    SS7[19][29] = 4'hD;
    SS7[20][29] = 4'hD;
    SS7[21][29] = 4'hD;
    SS7[22][29] = 4'hD;
    SS7[23][29] = 4'hA;
    SS7[24][29] = 4'hA;
    SS7[25][29] = 4'hA;
    SS7[26][29] = 4'hC;
    SS7[27][29] = 4'hC;
    SS7[28][29] = 4'hC;
    SS7[29][29] = 4'hC;
    SS7[30][29] = 4'hC;
    SS7[31][29] = 4'hC;
    SS7[32][29] = 4'hC;
    SS7[33][29] = 4'h0;
    SS7[34][29] = 4'h0;
    SS7[35][29] = 4'h0;
    SS7[36][29] = 4'h0;
    SS7[37][29] = 4'h0;
    SS7[38][29] = 4'h0;
    SS7[39][29] = 4'h0;
    SS7[40][29] = 4'h0;
    SS7[41][29] = 4'h0;
    SS7[42][29] = 4'h0;
    SS7[43][29] = 4'h0;
    SS7[44][29] = 4'h0;
    SS7[45][29] = 4'h0;
    SS7[46][29] = 4'h0;
    SS7[47][29] = 4'h0;
    SS7[0][30] = 4'h0;
    SS7[1][30] = 4'h0;
    SS7[2][30] = 4'h0;
    SS7[3][30] = 4'h0;
    SS7[4][30] = 4'h0;
    SS7[5][30] = 4'h0;
    SS7[6][30] = 4'h0;
    SS7[7][30] = 4'h3;
    SS7[8][30] = 4'h0;
    SS7[9][30] = 4'h0;
    SS7[10][30] = 4'h0;
    SS7[11][30] = 4'h0;
    SS7[12][30] = 4'h0;
    SS7[13][30] = 4'h0;
    SS7[14][30] = 4'hD;
    SS7[15][30] = 4'hD;
    SS7[16][30] = 4'h3;
    SS7[17][30] = 4'hD;
    SS7[18][30] = 4'hD;
    SS7[19][30] = 4'hD;
    SS7[20][30] = 4'hD;
    SS7[21][30] = 4'hD;
    SS7[22][30] = 4'hD;
    SS7[23][30] = 4'hA;
    SS7[24][30] = 4'hC;
    SS7[25][30] = 4'hC;
    SS7[26][30] = 4'hC;
    SS7[27][30] = 4'hC;
    SS7[28][30] = 4'hC;
    SS7[29][30] = 4'hC;
    SS7[30][30] = 4'hC;
    SS7[31][30] = 4'hC;
    SS7[32][30] = 4'hD;
    SS7[33][30] = 4'h0;
    SS7[34][30] = 4'h0;
    SS7[35][30] = 4'h0;
    SS7[36][30] = 4'h0;
    SS7[37][30] = 4'h0;
    SS7[38][30] = 4'h0;
    SS7[39][30] = 4'h0;
    SS7[40][30] = 4'h0;
    SS7[41][30] = 4'h0;
    SS7[42][30] = 4'h0;
    SS7[43][30] = 4'h0;
    SS7[44][30] = 4'h0;
    SS7[45][30] = 4'h0;
    SS7[46][30] = 4'h0;
    SS7[47][30] = 4'h0;
    SS7[0][31] = 4'h0;
    SS7[1][31] = 4'h0;
    SS7[2][31] = 4'h0;
    SS7[3][31] = 4'h0;
    SS7[4][31] = 4'h0;
    SS7[5][31] = 4'h0;
    SS7[6][31] = 4'h0;
    SS7[7][31] = 4'h0;
    SS7[8][31] = 4'h0;
    SS7[9][31] = 4'h0;
    SS7[10][31] = 4'h0;
    SS7[11][31] = 4'h0;
    SS7[12][31] = 4'h0;
    SS7[13][31] = 4'h0;
    SS7[14][31] = 4'h3;
    SS7[15][31] = 4'h3;
    SS7[16][31] = 4'h3;
    SS7[17][31] = 4'hD;
    SS7[18][31] = 4'hD;
    SS7[19][31] = 4'hD;
    SS7[20][31] = 4'hD;
    SS7[21][31] = 4'hC;
    SS7[22][31] = 4'hC;
    SS7[23][31] = 4'hC;
    SS7[24][31] = 4'hC;
    SS7[25][31] = 4'hC;
    SS7[26][31] = 4'hC;
    SS7[27][31] = 4'hC;
    SS7[28][31] = 4'hC;
    SS7[29][31] = 4'hC;
    SS7[30][31] = 4'hD;
    SS7[31][31] = 4'hD;
    SS7[32][31] = 4'hD;
    SS7[33][31] = 4'hD;
    SS7[34][31] = 4'h0;
    SS7[35][31] = 4'h0;
    SS7[36][31] = 4'h0;
    SS7[37][31] = 4'h0;
    SS7[38][31] = 4'h0;
    SS7[39][31] = 4'h0;
    SS7[40][31] = 4'h0;
    SS7[41][31] = 4'h0;
    SS7[42][31] = 4'h0;
    SS7[43][31] = 4'h0;
    SS7[44][31] = 4'h0;
    SS7[45][31] = 4'h0;
    SS7[46][31] = 4'h0;
    SS7[47][31] = 4'h0;
    SS7[0][32] = 4'h0;
    SS7[1][32] = 4'h0;
    SS7[2][32] = 4'h0;
    SS7[3][32] = 4'h0;
    SS7[4][32] = 4'h0;
    SS7[5][32] = 4'h0;
    SS7[6][32] = 4'h0;
    SS7[7][32] = 4'h0;
    SS7[8][32] = 4'h0;
    SS7[9][32] = 4'h0;
    SS7[10][32] = 4'h0;
    SS7[11][32] = 4'h0;
    SS7[12][32] = 4'h0;
    SS7[13][32] = 4'h0;
    SS7[14][32] = 4'h0;
    SS7[15][32] = 4'h3;
    SS7[16][32] = 4'h3;
    SS7[17][32] = 4'h3;
    SS7[18][32] = 4'hD;
    SS7[19][32] = 4'h0;
    SS7[20][32] = 4'h0;
    SS7[21][32] = 4'hC;
    SS7[22][32] = 4'hC;
    SS7[23][32] = 4'hC;
    SS7[24][32] = 4'hC;
    SS7[25][32] = 4'hC;
    SS7[26][32] = 4'hC;
    SS7[27][32] = 4'hC;
    SS7[28][32] = 4'hC;
    SS7[29][32] = 4'hC;
    SS7[30][32] = 4'hC;
    SS7[31][32] = 4'hD;
    SS7[32][32] = 4'hD;
    SS7[33][32] = 4'hD;
    SS7[34][32] = 4'h0;
    SS7[35][32] = 4'h0;
    SS7[36][32] = 4'h0;
    SS7[37][32] = 4'h0;
    SS7[38][32] = 4'h0;
    SS7[39][32] = 4'h0;
    SS7[40][32] = 4'h0;
    SS7[41][32] = 4'h0;
    SS7[42][32] = 4'h0;
    SS7[43][32] = 4'h0;
    SS7[44][32] = 4'h0;
    SS7[45][32] = 4'h0;
    SS7[46][32] = 4'h0;
    SS7[47][32] = 4'h0;
    SS7[0][33] = 4'h0;
    SS7[1][33] = 4'h0;
    SS7[2][33] = 4'h0;
    SS7[3][33] = 4'h0;
    SS7[4][33] = 4'h0;
    SS7[5][33] = 4'h0;
    SS7[6][33] = 4'h0;
    SS7[7][33] = 4'h0;
    SS7[8][33] = 4'h0;
    SS7[9][33] = 4'h0;
    SS7[10][33] = 4'h0;
    SS7[11][33] = 4'h0;
    SS7[12][33] = 4'h0;
    SS7[13][33] = 4'h0;
    SS7[14][33] = 4'h0;
    SS7[15][33] = 4'h3;
    SS7[16][33] = 4'h3;
    SS7[17][33] = 4'h0;
    SS7[18][33] = 4'h0;
    SS7[19][33] = 4'h0;
    SS7[20][33] = 4'h0;
    SS7[21][33] = 4'hE;
    SS7[22][33] = 4'hC;
    SS7[23][33] = 4'hC;
    SS7[24][33] = 4'hD;
    SS7[25][33] = 4'hC;
    SS7[26][33] = 4'hC;
    SS7[27][33] = 4'hC;
    SS7[28][33] = 4'hC;
    SS7[29][33] = 4'hC;
    SS7[30][33] = 4'hC;
    SS7[31][33] = 4'hD;
    SS7[32][33] = 4'hD;
    SS7[33][33] = 4'hD;
    SS7[34][33] = 4'h0;
    SS7[35][33] = 4'h0;
    SS7[36][33] = 4'h0;
    SS7[37][33] = 4'h0;
    SS7[38][33] = 4'h0;
    SS7[39][33] = 4'h0;
    SS7[40][33] = 4'h0;
    SS7[41][33] = 4'h0;
    SS7[42][33] = 4'h0;
    SS7[43][33] = 4'h0;
    SS7[44][33] = 4'h0;
    SS7[45][33] = 4'h0;
    SS7[46][33] = 4'h0;
    SS7[47][33] = 4'h0;
    SS7[0][34] = 4'h0;
    SS7[1][34] = 4'h0;
    SS7[2][34] = 4'h0;
    SS7[3][34] = 4'h0;
    SS7[4][34] = 4'h0;
    SS7[5][34] = 4'h0;
    SS7[6][34] = 4'h0;
    SS7[7][34] = 4'h0;
    SS7[8][34] = 4'h0;
    SS7[9][34] = 4'h0;
    SS7[10][34] = 4'h0;
    SS7[11][34] = 4'h0;
    SS7[12][34] = 4'h0;
    SS7[13][34] = 4'h0;
    SS7[14][34] = 4'h0;
    SS7[15][34] = 4'h0;
    SS7[16][34] = 4'h0;
    SS7[17][34] = 4'h0;
    SS7[18][34] = 4'h0;
    SS7[19][34] = 4'h0;
    SS7[20][34] = 4'h0;
    SS7[21][34] = 4'h0;
    SS7[22][34] = 4'hD;
    SS7[23][34] = 4'hD;
    SS7[24][34] = 4'hD;
    SS7[25][34] = 4'hC;
    SS7[26][34] = 4'hC;
    SS7[27][34] = 4'hC;
    SS7[28][34] = 4'hC;
    SS7[29][34] = 4'hC;
    SS7[30][34] = 4'hC;
    SS7[31][34] = 4'hC;
    SS7[32][34] = 4'hD;
    SS7[33][34] = 4'hD;
    SS7[34][34] = 4'hD;
    SS7[35][34] = 4'h0;
    SS7[36][34] = 4'h0;
    SS7[37][34] = 4'h0;
    SS7[38][34] = 4'h0;
    SS7[39][34] = 4'h0;
    SS7[40][34] = 4'h0;
    SS7[41][34] = 4'h0;
    SS7[42][34] = 4'h0;
    SS7[43][34] = 4'h0;
    SS7[44][34] = 4'h0;
    SS7[45][34] = 4'h0;
    SS7[46][34] = 4'h0;
    SS7[47][34] = 4'h0;
    SS7[0][35] = 4'h0;
    SS7[1][35] = 4'h0;
    SS7[2][35] = 4'h0;
    SS7[3][35] = 4'h0;
    SS7[4][35] = 4'h0;
    SS7[5][35] = 4'h0;
    SS7[6][35] = 4'h0;
    SS7[7][35] = 4'h0;
    SS7[8][35] = 4'h0;
    SS7[9][35] = 4'h0;
    SS7[10][35] = 4'h0;
    SS7[11][35] = 4'h0;
    SS7[12][35] = 4'h0;
    SS7[13][35] = 4'h0;
    SS7[14][35] = 4'h0;
    SS7[15][35] = 4'h0;
    SS7[16][35] = 4'h0;
    SS7[17][35] = 4'h0;
    SS7[18][35] = 4'h0;
    SS7[19][35] = 4'h0;
    SS7[20][35] = 4'h0;
    SS7[21][35] = 4'h0;
    SS7[22][35] = 4'hD;
    SS7[23][35] = 4'hD;
    SS7[24][35] = 4'hD;
    SS7[25][35] = 4'hD;
    SS7[26][35] = 4'hC;
    SS7[27][35] = 4'hC;
    SS7[28][35] = 4'hC;
    SS7[29][35] = 4'hC;
    SS7[30][35] = 4'hC;
    SS7[31][35] = 4'hC;
    SS7[32][35] = 4'hD;
    SS7[33][35] = 4'hD;
    SS7[34][35] = 4'hD;
    SS7[35][35] = 4'h0;
    SS7[36][35] = 4'h0;
    SS7[37][35] = 4'h0;
    SS7[38][35] = 4'h0;
    SS7[39][35] = 4'h0;
    SS7[40][35] = 4'h0;
    SS7[41][35] = 4'h0;
    SS7[42][35] = 4'h0;
    SS7[43][35] = 4'h0;
    SS7[44][35] = 4'h0;
    SS7[45][35] = 4'h0;
    SS7[46][35] = 4'h0;
    SS7[47][35] = 4'h0;
    SS7[0][36] = 4'h0;
    SS7[1][36] = 4'h0;
    SS7[2][36] = 4'h0;
    SS7[3][36] = 4'h0;
    SS7[4][36] = 4'h0;
    SS7[5][36] = 4'h0;
    SS7[6][36] = 4'h0;
    SS7[7][36] = 4'h0;
    SS7[8][36] = 4'h0;
    SS7[9][36] = 4'h0;
    SS7[10][36] = 4'h0;
    SS7[11][36] = 4'h0;
    SS7[12][36] = 4'h0;
    SS7[13][36] = 4'h0;
    SS7[14][36] = 4'h0;
    SS7[15][36] = 4'h0;
    SS7[16][36] = 4'h0;
    SS7[17][36] = 4'h0;
    SS7[18][36] = 4'h0;
    SS7[19][36] = 4'h0;
    SS7[20][36] = 4'h0;
    SS7[21][36] = 4'h0;
    SS7[22][36] = 4'h0;
    SS7[23][36] = 4'hD;
    SS7[24][36] = 4'hD;
    SS7[25][36] = 4'hD;
    SS7[26][36] = 4'hC;
    SS7[27][36] = 4'hC;
    SS7[28][36] = 4'hC;
    SS7[29][36] = 4'hC;
    SS7[30][36] = 4'hC;
    SS7[31][36] = 4'hC;
    SS7[32][36] = 4'hD;
    SS7[33][36] = 4'hD;
    SS7[34][36] = 4'hD;
    SS7[35][36] = 4'hD;
    SS7[36][36] = 4'h0;
    SS7[37][36] = 4'h0;
    SS7[38][36] = 4'h0;
    SS7[39][36] = 4'h0;
    SS7[40][36] = 4'h0;
    SS7[41][36] = 4'h0;
    SS7[42][36] = 4'h0;
    SS7[43][36] = 4'h0;
    SS7[44][36] = 4'h0;
    SS7[45][36] = 4'h0;
    SS7[46][36] = 4'h0;
    SS7[47][36] = 4'h0;
    SS7[0][37] = 4'h0;
    SS7[1][37] = 4'h0;
    SS7[2][37] = 4'h0;
    SS7[3][37] = 4'h0;
    SS7[4][37] = 4'h0;
    SS7[5][37] = 4'h0;
    SS7[6][37] = 4'h0;
    SS7[7][37] = 4'h0;
    SS7[8][37] = 4'h0;
    SS7[9][37] = 4'h0;
    SS7[10][37] = 4'h0;
    SS7[11][37] = 4'h0;
    SS7[12][37] = 4'h0;
    SS7[13][37] = 4'h0;
    SS7[14][37] = 4'h0;
    SS7[15][37] = 4'h0;
    SS7[16][37] = 4'h0;
    SS7[17][37] = 4'h0;
    SS7[18][37] = 4'h0;
    SS7[19][37] = 4'h0;
    SS7[20][37] = 4'h0;
    SS7[21][37] = 4'h0;
    SS7[22][37] = 4'h0;
    SS7[23][37] = 4'hD;
    SS7[24][37] = 4'hD;
    SS7[25][37] = 4'hD;
    SS7[26][37] = 4'hC;
    SS7[27][37] = 4'hC;
    SS7[28][37] = 4'hC;
    SS7[29][37] = 4'hC;
    SS7[30][37] = 4'hC;
    SS7[31][37] = 4'hC;
    SS7[32][37] = 4'hC;
    SS7[33][37] = 4'hD;
    SS7[34][37] = 4'hD;
    SS7[35][37] = 4'hD;
    SS7[36][37] = 4'h0;
    SS7[37][37] = 4'h0;
    SS7[38][37] = 4'h0;
    SS7[39][37] = 4'h0;
    SS7[40][37] = 4'h0;
    SS7[41][37] = 4'h0;
    SS7[42][37] = 4'h0;
    SS7[43][37] = 4'h0;
    SS7[44][37] = 4'h0;
    SS7[45][37] = 4'h0;
    SS7[46][37] = 4'h0;
    SS7[47][37] = 4'h0;
    SS7[0][38] = 4'h0;
    SS7[1][38] = 4'h0;
    SS7[2][38] = 4'h0;
    SS7[3][38] = 4'h0;
    SS7[4][38] = 4'h0;
    SS7[5][38] = 4'h0;
    SS7[6][38] = 4'h0;
    SS7[7][38] = 4'h0;
    SS7[8][38] = 4'h0;
    SS7[9][38] = 4'h0;
    SS7[10][38] = 4'h0;
    SS7[11][38] = 4'h0;
    SS7[12][38] = 4'h0;
    SS7[13][38] = 4'h0;
    SS7[14][38] = 4'h0;
    SS7[15][38] = 4'h0;
    SS7[16][38] = 4'h0;
    SS7[17][38] = 4'h0;
    SS7[18][38] = 4'h0;
    SS7[19][38] = 4'h0;
    SS7[20][38] = 4'h0;
    SS7[21][38] = 4'h0;
    SS7[22][38] = 4'h0;
    SS7[23][38] = 4'h0;
    SS7[24][38] = 4'hD;
    SS7[25][38] = 4'hD;
    SS7[26][38] = 4'hD;
    SS7[27][38] = 4'hC;
    SS7[28][38] = 4'hC;
    SS7[29][38] = 4'hC;
    SS7[30][38] = 4'hC;
    SS7[31][38] = 4'hC;
    SS7[32][38] = 4'hC;
    SS7[33][38] = 4'hD;
    SS7[34][38] = 4'hD;
    SS7[35][38] = 4'hF;
    SS7[36][38] = 4'h0;
    SS7[37][38] = 4'h0;
    SS7[38][38] = 4'h0;
    SS7[39][38] = 4'h0;
    SS7[40][38] = 4'h0;
    SS7[41][38] = 4'h0;
    SS7[42][38] = 4'h0;
    SS7[43][38] = 4'h0;
    SS7[44][38] = 4'h0;
    SS7[45][38] = 4'h0;
    SS7[46][38] = 4'h0;
    SS7[47][38] = 4'h0;
    SS7[0][39] = 4'h0;
    SS7[1][39] = 4'h0;
    SS7[2][39] = 4'h0;
    SS7[3][39] = 4'h0;
    SS7[4][39] = 4'h0;
    SS7[5][39] = 4'h0;
    SS7[6][39] = 4'h0;
    SS7[7][39] = 4'h0;
    SS7[8][39] = 4'h0;
    SS7[9][39] = 4'h0;
    SS7[10][39] = 4'h0;
    SS7[11][39] = 4'h0;
    SS7[12][39] = 4'h0;
    SS7[13][39] = 4'h0;
    SS7[14][39] = 4'h0;
    SS7[15][39] = 4'h0;
    SS7[16][39] = 4'h0;
    SS7[17][39] = 4'h0;
    SS7[18][39] = 4'h0;
    SS7[19][39] = 4'h0;
    SS7[20][39] = 4'h0;
    SS7[21][39] = 4'h0;
    SS7[22][39] = 4'h0;
    SS7[23][39] = 4'h0;
    SS7[24][39] = 4'hD;
    SS7[25][39] = 4'hD;
    SS7[26][39] = 4'hD;
    SS7[27][39] = 4'hC;
    SS7[28][39] = 4'hC;
    SS7[29][39] = 4'hC;
    SS7[30][39] = 4'hC;
    SS7[31][39] = 4'hC;
    SS7[32][39] = 4'hC;
    SS7[33][39] = 4'hC;
    SS7[34][39] = 4'h0;
    SS7[35][39] = 4'h0;
    SS7[36][39] = 4'h0;
    SS7[37][39] = 4'h0;
    SS7[38][39] = 4'h0;
    SS7[39][39] = 4'h0;
    SS7[40][39] = 4'h0;
    SS7[41][39] = 4'h0;
    SS7[42][39] = 4'h0;
    SS7[43][39] = 4'h0;
    SS7[44][39] = 4'h0;
    SS7[45][39] = 4'h0;
    SS7[46][39] = 4'h0;
    SS7[47][39] = 4'h0;
    SS7[0][40] = 4'h0;
    SS7[1][40] = 4'h0;
    SS7[2][40] = 4'h0;
    SS7[3][40] = 4'h0;
    SS7[4][40] = 4'h0;
    SS7[5][40] = 4'h0;
    SS7[6][40] = 4'h0;
    SS7[7][40] = 4'h0;
    SS7[8][40] = 4'h0;
    SS7[9][40] = 4'h0;
    SS7[10][40] = 4'h0;
    SS7[11][40] = 4'h0;
    SS7[12][40] = 4'h0;
    SS7[13][40] = 4'h0;
    SS7[14][40] = 4'h0;
    SS7[15][40] = 4'h0;
    SS7[16][40] = 4'h0;
    SS7[17][40] = 4'h0;
    SS7[18][40] = 4'h0;
    SS7[19][40] = 4'h0;
    SS7[20][40] = 4'h0;
    SS7[21][40] = 4'h0;
    SS7[22][40] = 4'h0;
    SS7[23][40] = 4'h0;
    SS7[24][40] = 4'hD;
    SS7[25][40] = 4'hD;
    SS7[26][40] = 4'hD;
    SS7[27][40] = 4'hD;
    SS7[28][40] = 4'hC;
    SS7[29][40] = 4'hC;
    SS7[30][40] = 4'hC;
    SS7[31][40] = 4'hC;
    SS7[32][40] = 4'hC;
    SS7[33][40] = 4'hC;
    SS7[34][40] = 4'h0;
    SS7[35][40] = 4'h0;
    SS7[36][40] = 4'h0;
    SS7[37][40] = 4'h0;
    SS7[38][40] = 4'h0;
    SS7[39][40] = 4'h0;
    SS7[40][40] = 4'h0;
    SS7[41][40] = 4'h0;
    SS7[42][40] = 4'h0;
    SS7[43][40] = 4'h0;
    SS7[44][40] = 4'h0;
    SS7[45][40] = 4'h0;
    SS7[46][40] = 4'h0;
    SS7[47][40] = 4'h0;
    SS7[0][41] = 4'h0;
    SS7[1][41] = 4'h0;
    SS7[2][41] = 4'h0;
    SS7[3][41] = 4'h0;
    SS7[4][41] = 4'h0;
    SS7[5][41] = 4'h0;
    SS7[6][41] = 4'h0;
    SS7[7][41] = 4'h0;
    SS7[8][41] = 4'h0;
    SS7[9][41] = 4'h0;
    SS7[10][41] = 4'h0;
    SS7[11][41] = 4'h0;
    SS7[12][41] = 4'h0;
    SS7[13][41] = 4'h0;
    SS7[14][41] = 4'h0;
    SS7[15][41] = 4'h0;
    SS7[16][41] = 4'h0;
    SS7[17][41] = 4'h0;
    SS7[18][41] = 4'h0;
    SS7[19][41] = 4'h0;
    SS7[20][41] = 4'h0;
    SS7[21][41] = 4'h0;
    SS7[22][41] = 4'h0;
    SS7[23][41] = 4'h0;
    SS7[24][41] = 4'h0;
    SS7[25][41] = 4'hD;
    SS7[26][41] = 4'hD;
    SS7[27][41] = 4'hD;
    SS7[28][41] = 4'hC;
    SS7[29][41] = 4'hC;
    SS7[30][41] = 4'hC;
    SS7[31][41] = 4'hC;
    SS7[32][41] = 4'hC;
    SS7[33][41] = 4'hC;
    SS7[34][41] = 4'h0;
    SS7[35][41] = 4'h0;
    SS7[36][41] = 4'h0;
    SS7[37][41] = 4'h0;
    SS7[38][41] = 4'h0;
    SS7[39][41] = 4'h0;
    SS7[40][41] = 4'h0;
    SS7[41][41] = 4'h0;
    SS7[42][41] = 4'h0;
    SS7[43][41] = 4'h0;
    SS7[44][41] = 4'h0;
    SS7[45][41] = 4'h0;
    SS7[46][41] = 4'h0;
    SS7[47][41] = 4'h0;
    SS7[0][42] = 4'h0;
    SS7[1][42] = 4'h0;
    SS7[2][42] = 4'h0;
    SS7[3][42] = 4'h0;
    SS7[4][42] = 4'h0;
    SS7[5][42] = 4'h0;
    SS7[6][42] = 4'h0;
    SS7[7][42] = 4'h0;
    SS7[8][42] = 4'h0;
    SS7[9][42] = 4'h0;
    SS7[10][42] = 4'h0;
    SS7[11][42] = 4'h0;
    SS7[12][42] = 4'h0;
    SS7[13][42] = 4'h0;
    SS7[14][42] = 4'h0;
    SS7[15][42] = 4'h0;
    SS7[16][42] = 4'h0;
    SS7[17][42] = 4'h0;
    SS7[18][42] = 4'h0;
    SS7[19][42] = 4'h0;
    SS7[20][42] = 4'h0;
    SS7[21][42] = 4'h0;
    SS7[22][42] = 4'h0;
    SS7[23][42] = 4'h0;
    SS7[24][42] = 4'h0;
    SS7[25][42] = 4'hD;
    SS7[26][42] = 4'h0;
    SS7[27][42] = 4'h0;
    SS7[28][42] = 4'hC;
    SS7[29][42] = 4'hC;
    SS7[30][42] = 4'hC;
    SS7[31][42] = 4'hC;
    SS7[32][42] = 4'hC;
    SS7[33][42] = 4'hC;
    SS7[34][42] = 4'hC;
    SS7[35][42] = 4'h0;
    SS7[36][42] = 4'h0;
    SS7[37][42] = 4'h0;
    SS7[38][42] = 4'h0;
    SS7[39][42] = 4'h0;
    SS7[40][42] = 4'h0;
    SS7[41][42] = 4'h0;
    SS7[42][42] = 4'h0;
    SS7[43][42] = 4'h0;
    SS7[44][42] = 4'h0;
    SS7[45][42] = 4'h0;
    SS7[46][42] = 4'h0;
    SS7[47][42] = 4'h0;
    SS7[0][43] = 4'h0;
    SS7[1][43] = 4'h0;
    SS7[2][43] = 4'h0;
    SS7[3][43] = 4'h0;
    SS7[4][43] = 4'h0;
    SS7[5][43] = 4'h0;
    SS7[6][43] = 4'h0;
    SS7[7][43] = 4'h0;
    SS7[8][43] = 4'h0;
    SS7[9][43] = 4'h0;
    SS7[10][43] = 4'h0;
    SS7[11][43] = 4'h0;
    SS7[12][43] = 4'h0;
    SS7[13][43] = 4'h0;
    SS7[14][43] = 4'h0;
    SS7[15][43] = 4'h0;
    SS7[16][43] = 4'h0;
    SS7[17][43] = 4'h0;
    SS7[18][43] = 4'h0;
    SS7[19][43] = 4'h0;
    SS7[20][43] = 4'h0;
    SS7[21][43] = 4'h0;
    SS7[22][43] = 4'h0;
    SS7[23][43] = 4'h0;
    SS7[24][43] = 4'h0;
    SS7[25][43] = 4'h0;
    SS7[26][43] = 4'h0;
    SS7[27][43] = 4'h0;
    SS7[28][43] = 4'h0;
    SS7[29][43] = 4'hC;
    SS7[30][43] = 4'hC;
    SS7[31][43] = 4'hC;
    SS7[32][43] = 4'hC;
    SS7[33][43] = 4'hC;
    SS7[34][43] = 4'hC;
    SS7[35][43] = 4'h0;
    SS7[36][43] = 4'h0;
    SS7[37][43] = 4'h0;
    SS7[38][43] = 4'h0;
    SS7[39][43] = 4'h0;
    SS7[40][43] = 4'h0;
    SS7[41][43] = 4'h0;
    SS7[42][43] = 4'h0;
    SS7[43][43] = 4'h0;
    SS7[44][43] = 4'h0;
    SS7[45][43] = 4'h0;
    SS7[46][43] = 4'h0;
    SS7[47][43] = 4'h0;
    SS7[0][44] = 4'h0;
    SS7[1][44] = 4'h0;
    SS7[2][44] = 4'h0;
    SS7[3][44] = 4'h0;
    SS7[4][44] = 4'h0;
    SS7[5][44] = 4'h0;
    SS7[6][44] = 4'h0;
    SS7[7][44] = 4'h0;
    SS7[8][44] = 4'h0;
    SS7[9][44] = 4'h0;
    SS7[10][44] = 4'h0;
    SS7[11][44] = 4'h0;
    SS7[12][44] = 4'h0;
    SS7[13][44] = 4'h0;
    SS7[14][44] = 4'h0;
    SS7[15][44] = 4'h0;
    SS7[16][44] = 4'h0;
    SS7[17][44] = 4'h0;
    SS7[18][44] = 4'h0;
    SS7[19][44] = 4'h0;
    SS7[20][44] = 4'h0;
    SS7[21][44] = 4'h0;
    SS7[22][44] = 4'h0;
    SS7[23][44] = 4'h0;
    SS7[24][44] = 4'h0;
    SS7[25][44] = 4'h0;
    SS7[26][44] = 4'h0;
    SS7[27][44] = 4'h0;
    SS7[28][44] = 4'h0;
    SS7[29][44] = 4'hC;
    SS7[30][44] = 4'hC;
    SS7[31][44] = 4'hC;
    SS7[32][44] = 4'hC;
    SS7[33][44] = 4'hC;
    SS7[34][44] = 4'hC;
    SS7[35][44] = 4'hC;
    SS7[36][44] = 4'h0;
    SS7[37][44] = 4'h0;
    SS7[38][44] = 4'h0;
    SS7[39][44] = 4'h0;
    SS7[40][44] = 4'h0;
    SS7[41][44] = 4'h0;
    SS7[42][44] = 4'h0;
    SS7[43][44] = 4'h0;
    SS7[44][44] = 4'h0;
    SS7[45][44] = 4'h0;
    SS7[46][44] = 4'h0;
    SS7[47][44] = 4'h0;
    SS7[0][45] = 4'h0;
    SS7[1][45] = 4'h0;
    SS7[2][45] = 4'h0;
    SS7[3][45] = 4'h0;
    SS7[4][45] = 4'h0;
    SS7[5][45] = 4'h0;
    SS7[6][45] = 4'h0;
    SS7[7][45] = 4'h0;
    SS7[8][45] = 4'h0;
    SS7[9][45] = 4'h0;
    SS7[10][45] = 4'h0;
    SS7[11][45] = 4'h0;
    SS7[12][45] = 4'h0;
    SS7[13][45] = 4'h0;
    SS7[14][45] = 4'h0;
    SS7[15][45] = 4'h0;
    SS7[16][45] = 4'h0;
    SS7[17][45] = 4'h0;
    SS7[18][45] = 4'h0;
    SS7[19][45] = 4'h0;
    SS7[20][45] = 4'h0;
    SS7[21][45] = 4'h0;
    SS7[22][45] = 4'h0;
    SS7[23][45] = 4'h0;
    SS7[24][45] = 4'h0;
    SS7[25][45] = 4'h0;
    SS7[26][45] = 4'h0;
    SS7[27][45] = 4'h0;
    SS7[28][45] = 4'h0;
    SS7[29][45] = 4'h0;
    SS7[30][45] = 4'hC;
    SS7[31][45] = 4'hC;
    SS7[32][45] = 4'hC;
    SS7[33][45] = 4'hC;
    SS7[34][45] = 4'h0;
    SS7[35][45] = 4'h0;
    SS7[36][45] = 4'h0;
    SS7[37][45] = 4'h0;
    SS7[38][45] = 4'h0;
    SS7[39][45] = 4'h0;
    SS7[40][45] = 4'h0;
    SS7[41][45] = 4'h0;
    SS7[42][45] = 4'h0;
    SS7[43][45] = 4'h0;
    SS7[44][45] = 4'h0;
    SS7[45][45] = 4'h0;
    SS7[46][45] = 4'h0;
    SS7[47][45] = 4'h0;
    SS7[0][46] = 4'h0;
    SS7[1][46] = 4'h0;
    SS7[2][46] = 4'h0;
    SS7[3][46] = 4'h0;
    SS7[4][46] = 4'h0;
    SS7[5][46] = 4'h0;
    SS7[6][46] = 4'h0;
    SS7[7][46] = 4'h0;
    SS7[8][46] = 4'h0;
    SS7[9][46] = 4'h0;
    SS7[10][46] = 4'h0;
    SS7[11][46] = 4'h0;
    SS7[12][46] = 4'h0;
    SS7[13][46] = 4'h0;
    SS7[14][46] = 4'h0;
    SS7[15][46] = 4'h0;
    SS7[16][46] = 4'h0;
    SS7[17][46] = 4'h0;
    SS7[18][46] = 4'h0;
    SS7[19][46] = 4'h0;
    SS7[20][46] = 4'h0;
    SS7[21][46] = 4'h0;
    SS7[22][46] = 4'h0;
    SS7[23][46] = 4'h0;
    SS7[24][46] = 4'h0;
    SS7[25][46] = 4'h0;
    SS7[26][46] = 4'h0;
    SS7[27][46] = 4'h0;
    SS7[28][46] = 4'h0;
    SS7[29][46] = 4'h0;
    SS7[30][46] = 4'hC;
    SS7[31][46] = 4'hC;
    SS7[32][46] = 4'h0;
    SS7[33][46] = 4'h0;
    SS7[34][46] = 4'h0;
    SS7[35][46] = 4'h0;
    SS7[36][46] = 4'h0;
    SS7[37][46] = 4'h0;
    SS7[38][46] = 4'h0;
    SS7[39][46] = 4'h0;
    SS7[40][46] = 4'h0;
    SS7[41][46] = 4'h0;
    SS7[42][46] = 4'h0;
    SS7[43][46] = 4'h0;
    SS7[44][46] = 4'h0;
    SS7[45][46] = 4'h0;
    SS7[46][46] = 4'h0;
    SS7[47][46] = 4'h0;
    SS7[0][47] = 4'h0;
    SS7[1][47] = 4'h0;
    SS7[2][47] = 4'h0;
    SS7[3][47] = 4'h0;
    SS7[4][47] = 4'h0;
    SS7[5][47] = 4'h0;
    SS7[6][47] = 4'h0;
    SS7[7][47] = 4'h0;
    SS7[8][47] = 4'h0;
    SS7[9][47] = 4'h0;
    SS7[10][47] = 4'h0;
    SS7[11][47] = 4'h0;
    SS7[12][47] = 4'h0;
    SS7[13][47] = 4'h0;
    SS7[14][47] = 4'h0;
    SS7[15][47] = 4'h0;
    SS7[16][47] = 4'h0;
    SS7[17][47] = 4'h0;
    SS7[18][47] = 4'h0;
    SS7[19][47] = 4'h0;
    SS7[20][47] = 4'h0;
    SS7[21][47] = 4'h0;
    SS7[22][47] = 4'h0;
    SS7[23][47] = 4'h0;
    SS7[24][47] = 4'h0;
    SS7[25][47] = 4'h0;
    SS7[26][47] = 4'h0;
    SS7[27][47] = 4'h0;
    SS7[28][47] = 4'h0;
    SS7[29][47] = 4'h0;
    SS7[30][47] = 4'h0;
    SS7[31][47] = 4'h0;
    SS7[32][47] = 4'h0;
    SS7[33][47] = 4'h0;
    SS7[34][47] = 4'h0;
    SS7[35][47] = 4'h0;
    SS7[36][47] = 4'h0;
    SS7[37][47] = 4'h0;
    SS7[38][47] = 4'h0;
    SS7[39][47] = 4'h0;
    SS7[40][47] = 4'h0;
    SS7[41][47] = 4'h0;
    SS7[42][47] = 4'h0;
    SS7[43][47] = 4'h0;
    SS7[44][47] = 4'h0;
    SS7[45][47] = 4'h0;
    SS7[46][47] = 4'h0;
    SS7[47][47] = 4'h0;
 
//SS 8
    SS8[0][0] = 4'h0;
    SS8[1][0] = 4'h0;
    SS8[2][0] = 4'h0;
    SS8[3][0] = 4'h0;
    SS8[4][0] = 4'h0;
    SS8[5][0] = 4'h0;
    SS8[6][0] = 4'h0;
    SS8[7][0] = 4'h0;
    SS8[8][0] = 4'h0;
    SS8[9][0] = 4'h0;
    SS8[10][0] = 4'h0;
    SS8[11][0] = 4'h0;
    SS8[12][0] = 4'h0;
    SS8[13][0] = 4'h0;
    SS8[14][0] = 4'h0;
    SS8[15][0] = 4'h0;
    SS8[16][0] = 4'h0;
    SS8[17][0] = 4'h0;
    SS8[18][0] = 4'h0;
    SS8[19][0] = 4'h0;
    SS8[20][0] = 4'h0;
    SS8[21][0] = 4'h0;
    SS8[22][0] = 4'h0;
    SS8[23][0] = 4'h0;
    SS8[24][0] = 4'h0;
    SS8[25][0] = 4'h0;
    SS8[26][0] = 4'hC;
    SS8[27][0] = 4'hC;
    SS8[28][0] = 4'hC;
    SS8[29][0] = 4'hC;
    SS8[30][0] = 4'hE;
    SS8[31][0] = 4'h0;
    SS8[32][0] = 4'h0;
    SS8[33][0] = 4'h0;
    SS8[34][0] = 4'h0;
    SS8[35][0] = 4'h0;
    SS8[36][0] = 4'h0;
    SS8[37][0] = 4'h0;
    SS8[38][0] = 4'h0;
    SS8[39][0] = 4'h0;
    SS8[40][0] = 4'h0;
    SS8[41][0] = 4'h0;
    SS8[42][0] = 4'h0;
    SS8[43][0] = 4'h0;
    SS8[44][0] = 4'h0;
    SS8[45][0] = 4'h0;
    SS8[46][0] = 4'h0;
    SS8[47][0] = 4'h0;
    SS8[0][1] = 4'h0;
    SS8[1][1] = 4'h0;
    SS8[2][1] = 4'h0;
    SS8[3][1] = 4'h0;
    SS8[4][1] = 4'h0;
    SS8[5][1] = 4'h0;
    SS8[6][1] = 4'h0;
    SS8[7][1] = 4'h0;
    SS8[8][1] = 4'h0;
    SS8[9][1] = 4'h0;
    SS8[10][1] = 4'h0;
    SS8[11][1] = 4'h0;
    SS8[12][1] = 4'h0;
    SS8[13][1] = 4'hD;
    SS8[14][1] = 4'h0;
    SS8[15][1] = 4'h0;
    SS8[16][1] = 4'h0;
    SS8[17][1] = 4'h0;
    SS8[18][1] = 4'h0;
    SS8[19][1] = 4'h0;
    SS8[20][1] = 4'h0;
    SS8[21][1] = 4'h0;
    SS8[22][1] = 4'h0;
    SS8[23][1] = 4'h0;
    SS8[24][1] = 4'h0;
    SS8[25][1] = 4'hC;
    SS8[26][1] = 4'hC;
    SS8[27][1] = 4'hC;
    SS8[28][1] = 4'hC;
    SS8[29][1] = 4'hC;
    SS8[30][1] = 4'hD;
    SS8[31][1] = 4'h0;
    SS8[32][1] = 4'h0;
    SS8[33][1] = 4'h0;
    SS8[34][1] = 4'h0;
    SS8[35][1] = 4'h0;
    SS8[36][1] = 4'h0;
    SS8[37][1] = 4'h0;
    SS8[38][1] = 4'h0;
    SS8[39][1] = 4'h0;
    SS8[40][1] = 4'h0;
    SS8[41][1] = 4'h0;
    SS8[42][1] = 4'h0;
    SS8[43][1] = 4'h0;
    SS8[44][1] = 4'h0;
    SS8[45][1] = 4'h0;
    SS8[46][1] = 4'h0;
    SS8[47][1] = 4'h0;
    SS8[0][2] = 4'h0;
    SS8[1][2] = 4'h0;
    SS8[2][2] = 4'h0;
    SS8[3][2] = 4'h0;
    SS8[4][2] = 4'h0;
    SS8[5][2] = 4'h0;
    SS8[6][2] = 4'h0;
    SS8[7][2] = 4'h0;
    SS8[8][2] = 4'h0;
    SS8[9][2] = 4'h0;
    SS8[10][2] = 4'h0;
    SS8[11][2] = 4'h0;
    SS8[12][2] = 4'hD;
    SS8[13][2] = 4'hD;
    SS8[14][2] = 4'hD;
    SS8[15][2] = 4'h0;
    SS8[16][2] = 4'h0;
    SS8[17][2] = 4'h0;
    SS8[18][2] = 4'h0;
    SS8[19][2] = 4'h0;
    SS8[20][2] = 4'h0;
    SS8[21][2] = 4'h0;
    SS8[22][2] = 4'h0;
    SS8[23][2] = 4'h0;
    SS8[24][2] = 4'hC;
    SS8[25][2] = 4'hC;
    SS8[26][2] = 4'hC;
    SS8[27][2] = 4'hC;
    SS8[28][2] = 4'hC;
    SS8[29][2] = 4'hD;
    SS8[30][2] = 4'hD;
    SS8[31][2] = 4'hD;
    SS8[32][2] = 4'h0;
    SS8[33][2] = 4'h0;
    SS8[34][2] = 4'h0;
    SS8[35][2] = 4'h0;
    SS8[36][2] = 4'h0;
    SS8[37][2] = 4'h0;
    SS8[38][2] = 4'h0;
    SS8[39][2] = 4'h0;
    SS8[40][2] = 4'h0;
    SS8[41][2] = 4'h0;
    SS8[42][2] = 4'h0;
    SS8[43][2] = 4'h0;
    SS8[44][2] = 4'h0;
    SS8[45][2] = 4'h0;
    SS8[46][2] = 4'h0;
    SS8[47][2] = 4'h0;
    SS8[0][3] = 4'h0;
    SS8[1][3] = 4'h0;
    SS8[2][3] = 4'h0;
    SS8[3][3] = 4'h0;
    SS8[4][3] = 4'h0;
    SS8[5][3] = 4'h0;
    SS8[6][3] = 4'h0;
    SS8[7][3] = 4'h0;
    SS8[8][3] = 4'h0;
    SS8[9][3] = 4'h0;
    SS8[10][3] = 4'h0;
    SS8[11][3] = 4'h0;
    SS8[12][3] = 4'hD;
    SS8[13][3] = 4'hD;
    SS8[14][3] = 4'hD;
    SS8[15][3] = 4'hD;
    SS8[16][3] = 4'h0;
    SS8[17][3] = 4'h0;
    SS8[18][3] = 4'h0;
    SS8[19][3] = 4'h0;
    SS8[20][3] = 4'h0;
    SS8[21][3] = 4'h0;
    SS8[22][3] = 4'h0;
    SS8[23][3] = 4'h0;
    SS8[24][3] = 4'h0;
    SS8[25][3] = 4'hC;
    SS8[26][3] = 4'hC;
    SS8[27][3] = 4'hC;
    SS8[28][3] = 4'hC;
    SS8[29][3] = 4'hD;
    SS8[30][3] = 4'hD;
    SS8[31][3] = 4'hD;
    SS8[32][3] = 4'h0;
    SS8[33][3] = 4'h0;
    SS8[34][3] = 4'h0;
    SS8[35][3] = 4'h0;
    SS8[36][3] = 4'h0;
    SS8[37][3] = 4'h0;
    SS8[38][3] = 4'h0;
    SS8[39][3] = 4'h0;
    SS8[40][3] = 4'h0;
    SS8[41][3] = 4'h0;
    SS8[42][3] = 4'h0;
    SS8[43][3] = 4'h0;
    SS8[44][3] = 4'h0;
    SS8[45][3] = 4'h0;
    SS8[46][3] = 4'h0;
    SS8[47][3] = 4'h0;
    SS8[0][4] = 4'h0;
    SS8[1][4] = 4'h0;
    SS8[2][4] = 4'h0;
    SS8[3][4] = 4'h0;
    SS8[4][4] = 4'h0;
    SS8[5][4] = 4'h0;
    SS8[6][4] = 4'h0;
    SS8[7][4] = 4'h0;
    SS8[8][4] = 4'h0;
    SS8[9][4] = 4'h0;
    SS8[10][4] = 4'h0;
    SS8[11][4] = 4'h0;
    SS8[12][4] = 4'h0;
    SS8[13][4] = 4'hD;
    SS8[14][4] = 4'hD;
    SS8[15][4] = 4'hD;
    SS8[16][4] = 4'hD;
    SS8[17][4] = 4'h0;
    SS8[18][4] = 4'h0;
    SS8[19][4] = 4'h0;
    SS8[20][4] = 4'h0;
    SS8[21][4] = 4'h0;
    SS8[22][4] = 4'h0;
    SS8[23][4] = 4'h0;
    SS8[24][4] = 4'h0;
    SS8[25][4] = 4'h0;
    SS8[26][4] = 4'hC;
    SS8[27][4] = 4'hC;
    SS8[28][4] = 4'hC;
    SS8[29][4] = 4'hC;
    SS8[30][4] = 4'hD;
    SS8[31][4] = 4'h0;
    SS8[32][4] = 4'h0;
    SS8[33][4] = 4'h0;
    SS8[34][4] = 4'h0;
    SS8[35][4] = 4'h0;
    SS8[36][4] = 4'h0;
    SS8[37][4] = 4'h0;
    SS8[38][4] = 4'h0;
    SS8[39][4] = 4'h0;
    SS8[40][4] = 4'h0;
    SS8[41][4] = 4'h0;
    SS8[42][4] = 4'h0;
    SS8[43][4] = 4'h0;
    SS8[44][4] = 4'h0;
    SS8[45][4] = 4'h0;
    SS8[46][4] = 4'h0;
    SS8[47][4] = 4'h0;
    SS8[0][5] = 4'h0;
    SS8[1][5] = 4'h0;
    SS8[2][5] = 4'h0;
    SS8[3][5] = 4'h0;
    SS8[4][5] = 4'h0;
    SS8[5][5] = 4'h0;
    SS8[6][5] = 4'h0;
    SS8[7][5] = 4'h0;
    SS8[8][5] = 4'h0;
    SS8[9][5] = 4'h0;
    SS8[10][5] = 4'h0;
    SS8[11][5] = 4'h0;
    SS8[12][5] = 4'h0;
    SS8[13][5] = 4'hD;
    SS8[14][5] = 4'hD;
    SS8[15][5] = 4'hD;
    SS8[16][5] = 4'hD;
    SS8[17][5] = 4'hE;
    SS8[18][5] = 4'h0;
    SS8[19][5] = 4'h0;
    SS8[20][5] = 4'h0;
    SS8[21][5] = 4'h0;
    SS8[22][5] = 4'h0;
    SS8[23][5] = 4'h0;
    SS8[24][5] = 4'h0;
    SS8[25][5] = 4'h0;
    SS8[26][5] = 4'hC;
    SS8[27][5] = 4'hC;
    SS8[28][5] = 4'hC;
    SS8[29][5] = 4'hC;
    SS8[30][5] = 4'hE;
    SS8[31][5] = 4'h0;
    SS8[32][5] = 4'h0;
    SS8[33][5] = 4'h0;
    SS8[34][5] = 4'h0;
    SS8[35][5] = 4'h0;
    SS8[36][5] = 4'h0;
    SS8[37][5] = 4'h0;
    SS8[38][5] = 4'h0;
    SS8[39][5] = 4'h0;
    SS8[40][5] = 4'h0;
    SS8[41][5] = 4'h0;
    SS8[42][5] = 4'h0;
    SS8[43][5] = 4'h0;
    SS8[44][5] = 4'h0;
    SS8[45][5] = 4'h0;
    SS8[46][5] = 4'h0;
    SS8[47][5] = 4'h0;
    SS8[0][6] = 4'h0;
    SS8[1][6] = 4'h0;
    SS8[2][6] = 4'h0;
    SS8[3][6] = 4'h0;
    SS8[4][6] = 4'h0;
    SS8[5][6] = 4'h0;
    SS8[6][6] = 4'h0;
    SS8[7][6] = 4'h0;
    SS8[8][6] = 4'h0;
    SS8[9][6] = 4'h0;
    SS8[10][6] = 4'h0;
    SS8[11][6] = 4'h0;
    SS8[12][6] = 4'hD;
    SS8[13][6] = 4'hD;
    SS8[14][6] = 4'hD;
    SS8[15][6] = 4'hD;
    SS8[16][6] = 4'hE;
    SS8[17][6] = 4'hE;
    SS8[18][6] = 4'hE;
    SS8[19][6] = 4'h0;
    SS8[20][6] = 4'h0;
    SS8[21][6] = 4'h0;
    SS8[22][6] = 4'h0;
    SS8[23][6] = 4'h0;
    SS8[24][6] = 4'h0;
    SS8[25][6] = 4'hC;
    SS8[26][6] = 4'hC;
    SS8[27][6] = 4'hC;
    SS8[28][6] = 4'hC;
    SS8[29][6] = 4'hE;
    SS8[30][6] = 4'hE;
    SS8[31][6] = 4'hE;
    SS8[32][6] = 4'h0;
    SS8[33][6] = 4'h0;
    SS8[34][6] = 4'h0;
    SS8[35][6] = 4'h0;
    SS8[36][6] = 4'h0;
    SS8[37][6] = 4'h0;
    SS8[38][6] = 4'h0;
    SS8[39][6] = 4'h0;
    SS8[40][6] = 4'h0;
    SS8[41][6] = 4'h0;
    SS8[42][6] = 4'h0;
    SS8[43][6] = 4'h0;
    SS8[44][6] = 4'h0;
    SS8[45][6] = 4'h0;
    SS8[46][6] = 4'h0;
    SS8[47][6] = 4'h0;
    SS8[0][7] = 4'h0;
    SS8[1][7] = 4'h0;
    SS8[2][7] = 4'h0;
    SS8[3][7] = 4'h0;
    SS8[4][7] = 4'h0;
    SS8[5][7] = 4'h0;
    SS8[6][7] = 4'h0;
    SS8[7][7] = 4'h0;
    SS8[8][7] = 4'h0;
    SS8[9][7] = 4'h0;
    SS8[10][7] = 4'h0;
    SS8[11][7] = 4'h0;
    SS8[12][7] = 4'hD;
    SS8[13][7] = 4'hD;
    SS8[14][7] = 4'hD;
    SS8[15][7] = 4'hD;
    SS8[16][7] = 4'hE;
    SS8[17][7] = 4'hE;
    SS8[18][7] = 4'hE;
    SS8[19][7] = 4'hE;
    SS8[20][7] = 4'h0;
    SS8[21][7] = 4'h0;
    SS8[22][7] = 4'h0;
    SS8[23][7] = 4'hD;
    SS8[24][7] = 4'hC;
    SS8[25][7] = 4'hC;
    SS8[26][7] = 4'hC;
    SS8[27][7] = 4'hC;
    SS8[28][7] = 4'hD;
    SS8[29][7] = 4'hE;
    SS8[30][7] = 4'hE;
    SS8[31][7] = 4'hE;
    SS8[32][7] = 4'h0;
    SS8[33][7] = 4'h0;
    SS8[34][7] = 4'h0;
    SS8[35][7] = 4'h0;
    SS8[36][7] = 4'h0;
    SS8[37][7] = 4'h0;
    SS8[38][7] = 4'h0;
    SS8[39][7] = 4'h0;
    SS8[40][7] = 4'h0;
    SS8[41][7] = 4'h0;
    SS8[42][7] = 4'h0;
    SS8[43][7] = 4'h0;
    SS8[44][7] = 4'h0;
    SS8[45][7] = 4'h0;
    SS8[46][7] = 4'h0;
    SS8[47][7] = 4'h0;
    SS8[0][8] = 4'h0;
    SS8[1][8] = 4'h0;
    SS8[2][8] = 4'h0;
    SS8[3][8] = 4'h0;
    SS8[4][8] = 4'h0;
    SS8[5][8] = 4'h0;
    SS8[6][8] = 4'h0;
    SS8[7][8] = 4'h0;
    SS8[8][8] = 4'h0;
    SS8[9][8] = 4'h0;
    SS8[10][8] = 4'h0;
    SS8[11][8] = 4'h0;
    SS8[12][8] = 4'h0;
    SS8[13][8] = 4'hD;
    SS8[14][8] = 4'hD;
    SS8[15][8] = 4'hD;
    SS8[16][8] = 4'hD;
    SS8[17][8] = 4'hE;
    SS8[18][8] = 4'hE;
    SS8[19][8] = 4'hE;
    SS8[20][8] = 4'hE;
    SS8[21][8] = 4'h0;
    SS8[22][8] = 4'hD;
    SS8[23][8] = 4'hC;
    SS8[24][8] = 4'hC;
    SS8[25][8] = 4'hC;
    SS8[26][8] = 4'hC;
    SS8[27][8] = 4'hD;
    SS8[28][8] = 4'hD;
    SS8[29][8] = 4'hD;
    SS8[30][8] = 4'hE;
    SS8[31][8] = 4'h0;
    SS8[32][8] = 4'h0;
    SS8[33][8] = 4'h0;
    SS8[34][8] = 4'h0;
    SS8[35][8] = 4'h0;
    SS8[36][8] = 4'h0;
    SS8[37][8] = 4'h0;
    SS8[38][8] = 4'h0;
    SS8[39][8] = 4'h0;
    SS8[40][8] = 4'h0;
    SS8[41][8] = 4'h0;
    SS8[42][8] = 4'h0;
    SS8[43][8] = 4'h0;
    SS8[44][8] = 4'h0;
    SS8[45][8] = 4'h0;
    SS8[46][8] = 4'h0;
    SS8[47][8] = 4'h0;
    SS8[0][9] = 4'h0;
    SS8[1][9] = 4'h0;
    SS8[2][9] = 4'h0;
    SS8[3][9] = 4'h0;
    SS8[4][9] = 4'h0;
    SS8[5][9] = 4'h0;
    SS8[6][9] = 4'h0;
    SS8[7][9] = 4'h0;
    SS8[8][9] = 4'h0;
    SS8[9][9] = 4'h0;
    SS8[10][9] = 4'h0;
    SS8[11][9] = 4'h0;
    SS8[12][9] = 4'h0;
    SS8[13][9] = 4'h3;
    SS8[14][9] = 4'hD;
    SS8[15][9] = 4'hD;
    SS8[16][9] = 4'hD;
    SS8[17][9] = 4'hE;
    SS8[18][9] = 4'hE;
    SS8[19][9] = 4'hE;
    SS8[20][9] = 4'hE;
    SS8[21][9] = 4'hE;
    SS8[22][9] = 4'hC;
    SS8[23][9] = 4'hC;
    SS8[24][9] = 4'hC;
    SS8[25][9] = 4'hC;
    SS8[26][9] = 4'hD;
    SS8[27][9] = 4'hD;
    SS8[28][9] = 4'hD;
    SS8[29][9] = 4'hD;
    SS8[30][9] = 4'hE;
    SS8[31][9] = 4'h0;
    SS8[32][9] = 4'h0;
    SS8[33][9] = 4'h0;
    SS8[34][9] = 4'h0;
    SS8[35][9] = 4'h0;
    SS8[36][9] = 4'h0;
    SS8[37][9] = 4'h0;
    SS8[38][9] = 4'h0;
    SS8[39][9] = 4'h0;
    SS8[40][9] = 4'h0;
    SS8[41][9] = 4'h0;
    SS8[42][9] = 4'h0;
    SS8[43][9] = 4'h0;
    SS8[44][9] = 4'h0;
    SS8[45][9] = 4'h0;
    SS8[46][9] = 4'h0;
    SS8[47][9] = 4'h0;
    SS8[0][10] = 4'h0;
    SS8[1][10] = 4'h0;
    SS8[2][10] = 4'h0;
    SS8[3][10] = 4'h0;
    SS8[4][10] = 4'h0;
    SS8[5][10] = 4'h0;
    SS8[6][10] = 4'h0;
    SS8[7][10] = 4'h0;
    SS8[8][10] = 4'h0;
    SS8[9][10] = 4'h0;
    SS8[10][10] = 4'h0;
    SS8[11][10] = 4'h0;
    SS8[12][10] = 4'h3;
    SS8[13][10] = 4'h3;
    SS8[14][10] = 4'h3;
    SS8[15][10] = 4'hD;
    SS8[16][10] = 4'hE;
    SS8[17][10] = 4'hE;
    SS8[18][10] = 4'hE;
    SS8[19][10] = 4'hE;
    SS8[20][10] = 4'hE;
    SS8[21][10] = 4'hC;
    SS8[22][10] = 4'hC;
    SS8[23][10] = 4'hC;
    SS8[24][10] = 4'hC;
    SS8[25][10] = 4'hC;
    SS8[26][10] = 4'hC;
    SS8[27][10] = 4'hD;
    SS8[28][10] = 4'hD;
    SS8[29][10] = 4'hE;
    SS8[30][10] = 4'hE;
    SS8[31][10] = 4'hE;
    SS8[32][10] = 4'h0;
    SS8[33][10] = 4'h0;
    SS8[34][10] = 4'h0;
    SS8[35][10] = 4'h0;
    SS8[36][10] = 4'h0;
    SS8[37][10] = 4'h0;
    SS8[38][10] = 4'h0;
    SS8[39][10] = 4'h0;
    SS8[40][10] = 4'h0;
    SS8[41][10] = 4'h0;
    SS8[42][10] = 4'h0;
    SS8[43][10] = 4'h0;
    SS8[44][10] = 4'h0;
    SS8[45][10] = 4'h0;
    SS8[46][10] = 4'h0;
    SS8[47][10] = 4'h0;
    SS8[0][11] = 4'h0;
    SS8[1][11] = 4'h0;
    SS8[2][11] = 4'h0;
    SS8[3][11] = 4'h0;
    SS8[4][11] = 4'h0;
    SS8[5][11] = 4'h0;
    SS8[6][11] = 4'h0;
    SS8[7][11] = 4'h0;
    SS8[8][11] = 4'h0;
    SS8[9][11] = 4'h0;
    SS8[10][11] = 4'h0;
    SS8[11][11] = 4'h2;
    SS8[12][11] = 4'h3;
    SS8[13][11] = 4'h3;
    SS8[14][11] = 4'h3;
    SS8[15][11] = 4'hD;
    SS8[16][11] = 4'hE;
    SS8[17][11] = 4'hE;
    SS8[18][11] = 4'hE;
    SS8[19][11] = 4'hE;
    SS8[20][11] = 4'hC;
    SS8[21][11] = 4'hC;
    SS8[22][11] = 4'hC;
    SS8[23][11] = 4'hC;
    SS8[24][11] = 4'hC;
    SS8[25][11] = 4'hC;
    SS8[26][11] = 4'hC;
    SS8[27][11] = 4'hC;
    SS8[28][11] = 4'hD;
    SS8[29][11] = 4'hE;
    SS8[30][11] = 4'hE;
    SS8[31][11] = 4'hE;
    SS8[32][11] = 4'h0;
    SS8[33][11] = 4'h0;
    SS8[34][11] = 4'h0;
    SS8[35][11] = 4'h0;
    SS8[36][11] = 4'h0;
    SS8[37][11] = 4'h0;
    SS8[38][11] = 4'h0;
    SS8[39][11] = 4'h0;
    SS8[40][11] = 4'h0;
    SS8[41][11] = 4'h0;
    SS8[42][11] = 4'h0;
    SS8[43][11] = 4'h0;
    SS8[44][11] = 4'h0;
    SS8[45][11] = 4'h0;
    SS8[46][11] = 4'h0;
    SS8[47][11] = 4'h0;
    SS8[0][12] = 4'h0;
    SS8[1][12] = 4'h0;
    SS8[2][12] = 4'h0;
    SS8[3][12] = 4'h0;
    SS8[4][12] = 4'h0;
    SS8[5][12] = 4'h0;
    SS8[6][12] = 4'h0;
    SS8[7][12] = 4'h0;
    SS8[8][12] = 4'h0;
    SS8[9][12] = 4'h0;
    SS8[10][12] = 4'h0;
    SS8[11][12] = 4'h0;
    SS8[12][12] = 4'h2;
    SS8[13][12] = 4'h3;
    SS8[14][12] = 4'hD;
    SS8[15][12] = 4'hD;
    SS8[16][12] = 4'hD;
    SS8[17][12] = 4'hE;
    SS8[18][12] = 4'hE;
    SS8[19][12] = 4'hE;
    SS8[20][12] = 4'hE;
    SS8[21][12] = 4'hC;
    SS8[22][12] = 4'hC;
    SS8[23][12] = 4'hC;
    SS8[24][12] = 4'hC;
    SS8[25][12] = 4'hC;
    SS8[26][12] = 4'hC;
    SS8[27][12] = 4'hD;
    SS8[28][12] = 4'hD;
    SS8[29][12] = 4'hD;
    SS8[30][12] = 4'hE;
    SS8[31][12] = 4'h0;
    SS8[32][12] = 4'h0;
    SS8[33][12] = 4'h0;
    SS8[34][12] = 4'h0;
    SS8[35][12] = 4'h0;
    SS8[36][12] = 4'h0;
    SS8[37][12] = 4'h0;
    SS8[38][12] = 4'h0;
    SS8[39][12] = 4'h0;
    SS8[40][12] = 4'h0;
    SS8[41][12] = 4'h0;
    SS8[42][12] = 4'h0;
    SS8[43][12] = 4'h0;
    SS8[44][12] = 4'h0;
    SS8[45][12] = 4'h0;
    SS8[46][12] = 4'h0;
    SS8[47][12] = 4'h0;
    SS8[0][13] = 4'h0;
    SS8[1][13] = 4'h0;
    SS8[2][13] = 4'h0;
    SS8[3][13] = 4'h0;
    SS8[4][13] = 4'h0;
    SS8[5][13] = 4'h0;
    SS8[6][13] = 4'h0;
    SS8[7][13] = 4'h0;
    SS8[8][13] = 4'h0;
    SS8[9][13] = 4'h0;
    SS8[10][13] = 4'h0;
    SS8[11][13] = 4'h0;
    SS8[12][13] = 4'h0;
    SS8[13][13] = 4'hE;
    SS8[14][13] = 4'hD;
    SS8[15][13] = 4'hD;
    SS8[16][13] = 4'hD;
    SS8[17][13] = 4'hD;
    SS8[18][13] = 4'hE;
    SS8[19][13] = 4'hE;
    SS8[20][13] = 4'hE;
    SS8[21][13] = 4'hE;
    SS8[22][13] = 4'hC;
    SS8[23][13] = 4'hC;
    SS8[24][13] = 4'hC;
    SS8[25][13] = 4'hC;
    SS8[26][13] = 4'hD;
    SS8[27][13] = 4'hD;
    SS8[28][13] = 4'hD;
    SS8[29][13] = 4'hD;
    SS8[30][13] = 4'h0;
    SS8[31][13] = 4'h0;
    SS8[32][13] = 4'h0;
    SS8[33][13] = 4'h0;
    SS8[34][13] = 4'h0;
    SS8[35][13] = 4'h0;
    SS8[36][13] = 4'h0;
    SS8[37][13] = 4'h0;
    SS8[38][13] = 4'h0;
    SS8[39][13] = 4'h0;
    SS8[40][13] = 4'h0;
    SS8[41][13] = 4'h0;
    SS8[42][13] = 4'h0;
    SS8[43][13] = 4'h0;
    SS8[44][13] = 4'h0;
    SS8[45][13] = 4'h0;
    SS8[46][13] = 4'h0;
    SS8[47][13] = 4'h0;
    SS8[0][14] = 4'h0;
    SS8[1][14] = 4'h0;
    SS8[2][14] = 4'h0;
    SS8[3][14] = 4'h0;
    SS8[4][14] = 4'h0;
    SS8[5][14] = 4'h0;
    SS8[6][14] = 4'h0;
    SS8[7][14] = 4'h0;
    SS8[8][14] = 4'h0;
    SS8[9][14] = 4'h0;
    SS8[10][14] = 4'h0;
    SS8[11][14] = 4'h0;
    SS8[12][14] = 4'h0;
    SS8[13][14] = 4'h0;
    SS8[14][14] = 4'hE;
    SS8[15][14] = 4'hD;
    SS8[16][14] = 4'hD;
    SS8[17][14] = 4'hD;
    SS8[18][14] = 4'hD;
    SS8[19][14] = 4'hE;
    SS8[20][14] = 4'hE;
    SS8[21][14] = 4'hC;
    SS8[22][14] = 4'hC;
    SS8[23][14] = 4'hC;
    SS8[24][14] = 4'hC;
    SS8[25][14] = 4'hC;
    SS8[26][14] = 4'hC;
    SS8[27][14] = 4'hD;
    SS8[28][14] = 4'hD;
    SS8[29][14] = 4'hE;
    SS8[30][14] = 4'hE;
    SS8[31][14] = 4'h0;
    SS8[32][14] = 4'h0;
    SS8[33][14] = 4'h0;
    SS8[34][14] = 4'h0;
    SS8[35][14] = 4'h0;
    SS8[36][14] = 4'h0;
    SS8[37][14] = 4'h0;
    SS8[38][14] = 4'h0;
    SS8[39][14] = 4'h0;
    SS8[40][14] = 4'h0;
    SS8[41][14] = 4'h0;
    SS8[42][14] = 4'h0;
    SS8[43][14] = 4'h0;
    SS8[44][14] = 4'h0;
    SS8[45][14] = 4'h0;
    SS8[46][14] = 4'h0;
    SS8[47][14] = 4'h0;
    SS8[0][15] = 4'h0;
    SS8[1][15] = 4'h0;
    SS8[2][15] = 4'h0;
    SS8[3][15] = 4'h0;
    SS8[4][15] = 4'h0;
    SS8[5][15] = 4'h0;
    SS8[6][15] = 4'h0;
    SS8[7][15] = 4'h0;
    SS8[8][15] = 4'h0;
    SS8[9][15] = 4'h0;
    SS8[10][15] = 4'h0;
    SS8[11][15] = 4'h0;
    SS8[12][15] = 4'h0;
    SS8[13][15] = 4'h0;
    SS8[14][15] = 4'h0;
    SS8[15][15] = 4'hD;
    SS8[16][15] = 4'hD;
    SS8[17][15] = 4'hD;
    SS8[18][15] = 4'hD;
    SS8[19][15] = 4'hD;
    SS8[20][15] = 4'hC;
    SS8[21][15] = 4'hC;
    SS8[22][15] = 4'hC;
    SS8[23][15] = 4'hC;
    SS8[24][15] = 4'hC;
    SS8[25][15] = 4'hC;
    SS8[26][15] = 4'hC;
    SS8[27][15] = 4'hC;
    SS8[28][15] = 4'hE;
    SS8[29][15] = 4'hE;
    SS8[30][15] = 4'hE;
    SS8[31][15] = 4'hE;
    SS8[32][15] = 4'hF;
    SS8[33][15] = 4'h0;
    SS8[34][15] = 4'h0;
    SS8[35][15] = 4'h0;
    SS8[36][15] = 4'h0;
    SS8[37][15] = 4'h0;
    SS8[38][15] = 4'h0;
    SS8[39][15] = 4'h0;
    SS8[40][15] = 4'h0;
    SS8[41][15] = 4'h0;
    SS8[42][15] = 4'h0;
    SS8[43][15] = 4'h0;
    SS8[44][15] = 4'h0;
    SS8[45][15] = 4'h0;
    SS8[46][15] = 4'h0;
    SS8[47][15] = 4'h0;
    SS8[0][16] = 4'h0;
    SS8[1][16] = 4'h0;
    SS8[2][16] = 4'h0;
    SS8[3][16] = 4'h0;
    SS8[4][16] = 4'h0;
    SS8[5][16] = 4'h0;
    SS8[6][16] = 4'h0;
    SS8[7][16] = 4'h0;
    SS8[8][16] = 4'h0;
    SS8[9][16] = 4'h0;
    SS8[10][16] = 4'h0;
    SS8[11][16] = 4'h0;
    SS8[12][16] = 4'h0;
    SS8[13][16] = 4'h0;
    SS8[14][16] = 4'h0;
    SS8[15][16] = 4'hD;
    SS8[16][16] = 4'hD;
    SS8[17][16] = 4'hD;
    SS8[18][16] = 4'hD;
    SS8[19][16] = 4'hE;
    SS8[20][16] = 4'hE;
    SS8[21][16] = 4'hC;
    SS8[22][16] = 4'hC;
    SS8[23][16] = 4'hC;
    SS8[24][16] = 4'hC;
    SS8[25][16] = 4'hC;
    SS8[26][16] = 4'hC;
    SS8[27][16] = 4'hE;
    SS8[28][16] = 4'hE;
    SS8[29][16] = 4'hE;
    SS8[30][16] = 4'hE;
    SS8[31][16] = 4'hE;
    SS8[32][16] = 4'hE;
    SS8[33][16] = 4'h0;
    SS8[34][16] = 4'h0;
    SS8[35][16] = 4'h0;
    SS8[36][16] = 4'hE;
    SS8[37][16] = 4'hE;
    SS8[38][16] = 4'h0;
    SS8[39][16] = 4'h0;
    SS8[40][16] = 4'hE;
    SS8[41][16] = 4'hE;
    SS8[42][16] = 4'h0;
    SS8[43][16] = 4'h0;
    SS8[44][16] = 4'hD;
    SS8[45][16] = 4'hD;
    SS8[46][16] = 4'h0;
    SS8[47][16] = 4'h0;
    SS8[0][17] = 4'h0;
    SS8[1][17] = 4'h0;
    SS8[2][17] = 4'h0;
    SS8[3][17] = 4'h0;
    SS8[4][17] = 4'h0;
    SS8[5][17] = 4'h0;
    SS8[6][17] = 4'h0;
    SS8[7][17] = 4'h0;
    SS8[8][17] = 4'h0;
    SS8[9][17] = 4'h0;
    SS8[10][17] = 4'h0;
    SS8[11][17] = 4'h0;
    SS8[12][17] = 4'h0;
    SS8[13][17] = 4'h0;
    SS8[14][17] = 4'hD;
    SS8[15][17] = 4'hD;
    SS8[16][17] = 4'hD;
    SS8[17][17] = 4'hD;
    SS8[18][17] = 4'hE;
    SS8[19][17] = 4'hE;
    SS8[20][17] = 4'hE;
    SS8[21][17] = 4'hE;
    SS8[22][17] = 4'hC;
    SS8[23][17] = 4'hC;
    SS8[24][17] = 4'hC;
    SS8[25][17] = 4'hC;
    SS8[26][17] = 4'hE;
    SS8[27][17] = 4'hE;
    SS8[28][17] = 4'hE;
    SS8[29][17] = 4'hE;
    SS8[30][17] = 4'hE;
    SS8[31][17] = 4'hE;
    SS8[32][17] = 4'hE;
    SS8[33][17] = 4'hE;
    SS8[34][17] = 4'h0;
    SS8[35][17] = 4'hE;
    SS8[36][17] = 4'hE;
    SS8[37][17] = 4'hE;
    SS8[38][17] = 4'hE;
    SS8[39][17] = 4'hE;
    SS8[40][17] = 4'hE;
    SS8[41][17] = 4'hE;
    SS8[42][17] = 4'hE;
    SS8[43][17] = 4'hD;
    SS8[44][17] = 4'hD;
    SS8[45][17] = 4'hD;
    SS8[46][17] = 4'hD;
    SS8[47][17] = 4'hE;
    SS8[0][18] = 4'h0;
    SS8[1][18] = 4'h0;
    SS8[2][18] = 4'h0;
    SS8[3][18] = 4'h0;
    SS8[4][18] = 4'h0;
    SS8[5][18] = 4'h0;
    SS8[6][18] = 4'h0;
    SS8[7][18] = 4'h0;
    SS8[8][18] = 4'h0;
    SS8[9][18] = 4'h0;
    SS8[10][18] = 4'h0;
    SS8[11][18] = 4'h0;
    SS8[12][18] = 4'h2;
    SS8[13][18] = 4'h3;
    SS8[14][18] = 4'hD;
    SS8[15][18] = 4'hD;
    SS8[16][18] = 4'hD;
    SS8[17][18] = 4'hD;
    SS8[18][18] = 4'hD;
    SS8[19][18] = 4'hE;
    SS8[20][18] = 4'hE;
    SS8[21][18] = 4'hC;
    SS8[22][18] = 4'hC;
    SS8[23][18] = 4'hC;
    SS8[24][18] = 4'hC;
    SS8[25][18] = 4'hD;
    SS8[26][18] = 4'hD;
    SS8[27][18] = 4'hE;
    SS8[28][18] = 4'hE;
    SS8[29][18] = 4'hE;
    SS8[30][18] = 4'hE;
    SS8[31][18] = 4'hE;
    SS8[32][18] = 4'hE;
    SS8[33][18] = 4'hE;
    SS8[34][18] = 4'hD;
    SS8[35][18] = 4'hD;
    SS8[36][18] = 4'hE;
    SS8[37][18] = 4'hE;
    SS8[38][18] = 4'hD;
    SS8[39][18] = 4'hD;
    SS8[40][18] = 4'hE;
    SS8[41][18] = 4'hE;
    SS8[42][18] = 4'hC;
    SS8[43][18] = 4'hC;
    SS8[44][18] = 4'hD;
    SS8[45][18] = 4'hD;
    SS8[46][18] = 4'hC;
    SS8[47][18] = 4'hC;
    SS8[0][19] = 4'h0;
    SS8[1][19] = 4'h0;
    SS8[2][19] = 4'h0;
    SS8[3][19] = 4'h0;
    SS8[4][19] = 4'h0;
    SS8[5][19] = 4'h0;
    SS8[6][19] = 4'h0;
    SS8[7][19] = 4'h0;
    SS8[8][19] = 4'h0;
    SS8[9][19] = 4'h0;
    SS8[10][19] = 4'h0;
    SS8[11][19] = 4'h2;
    SS8[12][19] = 4'h3;
    SS8[13][19] = 4'h3;
    SS8[14][19] = 4'h3;
    SS8[15][19] = 4'hD;
    SS8[16][19] = 4'hD;
    SS8[17][19] = 4'hD;
    SS8[18][19] = 4'hD;
    SS8[19][19] = 4'hD;
    SS8[20][19] = 4'hC;
    SS8[21][19] = 4'hC;
    SS8[22][19] = 4'hC;
    SS8[23][19] = 4'hC;
    SS8[24][19] = 4'hD;
    SS8[25][19] = 4'hD;
    SS8[26][19] = 4'hD;
    SS8[27][19] = 4'hD;
    SS8[28][19] = 4'hE;
    SS8[29][19] = 4'hE;
    SS8[30][19] = 4'hE;
    SS8[31][19] = 4'hE;
    SS8[32][19] = 4'hE;
    SS8[33][19] = 4'hD;
    SS8[34][19] = 4'hD;
    SS8[35][19] = 4'hD;
    SS8[36][19] = 4'hD;
    SS8[37][19] = 4'hD;
    SS8[38][19] = 4'hD;
    SS8[39][19] = 4'hD;
    SS8[40][19] = 4'hD;
    SS8[41][19] = 4'hC;
    SS8[42][19] = 4'hC;
    SS8[43][19] = 4'hC;
    SS8[44][19] = 4'hC;
    SS8[45][19] = 4'hC;
    SS8[46][19] = 4'hC;
    SS8[47][19] = 4'hC;
    SS8[0][20] = 4'h0;
    SS8[1][20] = 4'h0;
    SS8[2][20] = 4'h0;
    SS8[3][20] = 4'h0;
    SS8[4][20] = 4'h0;
    SS8[5][20] = 4'h0;
    SS8[6][20] = 4'h0;
    SS8[7][20] = 4'h0;
    SS8[8][20] = 4'h0;
    SS8[9][20] = 4'h0;
    SS8[10][20] = 4'h0;
    SS8[11][20] = 4'h0;
    SS8[12][20] = 4'h3;
    SS8[13][20] = 4'h3;
    SS8[14][20] = 4'h3;
    SS8[15][20] = 4'hD;
    SS8[16][20] = 4'hD;
    SS8[17][20] = 4'hD;
    SS8[18][20] = 4'hD;
    SS8[19][20] = 4'hC;
    SS8[20][20] = 4'hC;
    SS8[21][20] = 4'hC;
    SS8[22][20] = 4'hC;
    SS8[23][20] = 4'hC;
    SS8[24][20] = 4'hC;
    SS8[25][20] = 4'hD;
    SS8[26][20] = 4'hD;
    SS8[27][20] = 4'hD;
    SS8[28][20] = 4'hD;
    SS8[29][20] = 4'hE;
    SS8[30][20] = 4'hE;
    SS8[31][20] = 4'hE;
    SS8[32][20] = 4'hC;
    SS8[33][20] = 4'hD;
    SS8[34][20] = 4'hD;
    SS8[35][20] = 4'hD;
    SS8[36][20] = 4'hC;
    SS8[37][20] = 4'hD;
    SS8[38][20] = 4'hD;
    SS8[39][20] = 4'hD;
    SS8[40][20] = 4'hC;
    SS8[41][20] = 4'hC;
    SS8[42][20] = 4'hC;
    SS8[43][20] = 4'hC;
    SS8[44][20] = 4'hC;
    SS8[45][20] = 4'hC;
    SS8[46][20] = 4'hC;
    SS8[47][20] = 4'hC;
    SS8[0][21] = 4'h0;
    SS8[1][21] = 4'h0;
    SS8[2][21] = 4'h0;
    SS8[3][21] = 4'h0;
    SS8[4][21] = 4'h0;
    SS8[5][21] = 4'h0;
    SS8[6][21] = 4'h0;
    SS8[7][21] = 4'h0;
    SS8[8][21] = 4'h0;
    SS8[9][21] = 4'h0;
    SS8[10][21] = 4'h0;
    SS8[11][21] = 4'h0;
    SS8[12][21] = 4'h0;
    SS8[13][21] = 4'h3;
    SS8[14][21] = 4'hD;
    SS8[15][21] = 4'hD;
    SS8[16][21] = 4'hD;
    SS8[17][21] = 4'hD;
    SS8[18][21] = 4'hC;
    SS8[19][21] = 4'hC;
    SS8[20][21] = 4'hC;
    SS8[21][21] = 4'hC;
    SS8[22][21] = 4'hC;
    SS8[23][21] = 4'hC;
    SS8[24][21] = 4'hC;
    SS8[25][21] = 4'hC;
    SS8[26][21] = 4'hD;
    SS8[27][21] = 4'hD;
    SS8[28][21] = 4'hD;
    SS8[29][21] = 4'hD;
    SS8[30][21] = 4'hE;
    SS8[31][21] = 4'hC;
    SS8[32][21] = 4'hC;
    SS8[33][21] = 4'hC;
    SS8[34][21] = 4'hD;
    SS8[35][21] = 4'hC;
    SS8[36][21] = 4'hC;
    SS8[37][21] = 4'hC;
    SS8[38][21] = 4'hD;
    SS8[39][21] = 4'hC;
    SS8[40][21] = 4'hC;
    SS8[41][21] = 4'hC;
    SS8[42][21] = 4'hC;
    SS8[43][21] = 4'hC;
    SS8[44][21] = 4'hC;
    SS8[45][21] = 4'hC;
    SS8[46][21] = 4'hC;
    SS8[47][21] = 4'hC;
    SS8[0][22] = 4'h0;
    SS8[1][22] = 4'h0;
    SS8[2][22] = 4'h0;
    SS8[3][22] = 4'h0;
    SS8[4][22] = 4'h0;
    SS8[5][22] = 4'h0;
    SS8[6][22] = 4'h0;
    SS8[7][22] = 4'h0;
    SS8[8][22] = 4'h0;
    SS8[9][22] = 4'h0;
    SS8[10][22] = 4'h0;
    SS8[11][22] = 4'h0;
    SS8[12][22] = 4'h0;
    SS8[13][22] = 4'h0;
    SS8[14][22] = 4'hD;
    SS8[15][22] = 4'hD;
    SS8[16][22] = 4'hD;
    SS8[17][22] = 4'hD;
    SS8[18][22] = 4'hC;
    SS8[19][22] = 4'hC;
    SS8[20][22] = 4'hC;
    SS8[21][22] = 4'hD;
    SS8[22][22] = 4'hC;
    SS8[23][22] = 4'hC;
    SS8[24][22] = 4'hC;
    SS8[25][22] = 4'hC;
    SS8[26][22] = 4'hC;
    SS8[27][22] = 4'hD;
    SS8[28][22] = 4'hD;
    SS8[29][22] = 4'hD;
    SS8[30][22] = 4'hC;
    SS8[31][22] = 4'hC;
    SS8[32][22] = 4'hC;
    SS8[33][22] = 4'hC;
    SS8[34][22] = 4'hC;
    SS8[35][22] = 4'hC;
    SS8[36][22] = 4'hC;
    SS8[37][22] = 4'hC;
    SS8[38][22] = 4'hC;
    SS8[39][22] = 4'hC;
    SS8[40][22] = 4'hC;
    SS8[41][22] = 4'hC;
    SS8[42][22] = 4'h0;
    SS8[43][22] = 4'h0;
    SS8[44][22] = 4'hC;
    SS8[45][22] = 4'hC;
    SS8[46][22] = 4'hC;
    SS8[47][22] = 4'h0;
    SS8[0][23] = 4'h0;
    SS8[1][23] = 4'h0;
    SS8[2][23] = 4'h0;
    SS8[3][23] = 4'h0;
    SS8[4][23] = 4'h0;
    SS8[5][23] = 4'h0;
    SS8[6][23] = 4'h0;
    SS8[7][23] = 4'h0;
    SS8[8][23] = 4'h0;
    SS8[9][23] = 4'h0;
    SS8[10][23] = 4'h0;
    SS8[11][23] = 4'h0;
    SS8[12][23] = 4'h0;
    SS8[13][23] = 4'h0;
    SS8[14][23] = 4'h0;
    SS8[15][23] = 4'hD;
    SS8[16][23] = 4'hD;
    SS8[17][23] = 4'hD;
    SS8[18][23] = 4'hD;
    SS8[19][23] = 4'hC;
    SS8[20][23] = 4'hD;
    SS8[21][23] = 4'hD;
    SS8[22][23] = 4'hD;
    SS8[23][23] = 4'hC;
    SS8[24][23] = 4'hC;
    SS8[25][23] = 4'hC;
    SS8[26][23] = 4'hC;
    SS8[27][23] = 4'hC;
    SS8[28][23] = 4'hD;
    SS8[29][23] = 4'hC;
    SS8[30][23] = 4'hC;
    SS8[31][23] = 4'hC;
    SS8[32][23] = 4'hC;
    SS8[33][23] = 4'hC;
    SS8[34][23] = 4'hC;
    SS8[35][23] = 4'hC;
    SS8[36][23] = 4'hC;
    SS8[37][23] = 4'hC;
    SS8[38][23] = 4'hC;
    SS8[39][23] = 4'hC;
    SS8[40][23] = 4'hC;
    SS8[41][23] = 4'h0;
    SS8[42][23] = 4'h0;
    SS8[43][23] = 4'h0;
    SS8[44][23] = 4'h0;
    SS8[45][23] = 4'hC;
    SS8[46][23] = 4'h0;
    SS8[47][23] = 4'h0;
    SS8[0][24] = 4'h0;
    SS8[1][24] = 4'h0;
    SS8[2][24] = 4'h0;
    SS8[3][24] = 4'h0;
    SS8[4][24] = 4'h0;
    SS8[5][24] = 4'h0;
    SS8[6][24] = 4'h0;
    SS8[7][24] = 4'h0;
    SS8[8][24] = 4'h0;
    SS8[9][24] = 4'h0;
    SS8[10][24] = 4'h0;
    SS8[11][24] = 4'h0;
    SS8[12][24] = 4'h0;
    SS8[13][24] = 4'h0;
    SS8[14][24] = 4'h0;
    SS8[15][24] = 4'hC;
    SS8[16][24] = 4'hD;
    SS8[17][24] = 4'hD;
    SS8[18][24] = 4'hD;
    SS8[19][24] = 4'hA;
    SS8[20][24] = 4'hD;
    SS8[21][24] = 4'hD;
    SS8[22][24] = 4'hD;
    SS8[23][24] = 4'hD;
    SS8[24][24] = 4'hC;
    SS8[25][24] = 4'hC;
    SS8[26][24] = 4'hC;
    SS8[27][24] = 4'hC;
    SS8[28][24] = 4'hC;
    SS8[29][24] = 4'hC;
    SS8[30][24] = 4'hC;
    SS8[31][24] = 4'hC;
    SS8[32][24] = 4'hC;
    SS8[33][24] = 4'hC;
    SS8[34][24] = 4'hC;
    SS8[35][24] = 4'hC;
    SS8[36][24] = 4'hC;
    SS8[37][24] = 4'hC;
    SS8[38][24] = 4'hC;
    SS8[39][24] = 4'hC;
    SS8[40][24] = 4'hD;
    SS8[41][24] = 4'h0;
    SS8[42][24] = 4'h0;
    SS8[43][24] = 4'h0;
    SS8[44][24] = 4'h0;
    SS8[45][24] = 4'h0;
    SS8[46][24] = 4'h0;
    SS8[47][24] = 4'h0;
    SS8[0][25] = 4'h0;
    SS8[1][25] = 4'h0;
    SS8[2][25] = 4'h0;
    SS8[3][25] = 4'h0;
    SS8[4][25] = 4'h0;
    SS8[5][25] = 4'h0;
    SS8[6][25] = 4'h0;
    SS8[7][25] = 4'h0;
    SS8[8][25] = 4'h0;
    SS8[9][25] = 4'h0;
    SS8[10][25] = 4'h0;
    SS8[11][25] = 4'h0;
    SS8[12][25] = 4'h0;
    SS8[13][25] = 4'h0;
    SS8[14][25] = 4'hC;
    SS8[15][25] = 4'hC;
    SS8[16][25] = 4'hC;
    SS8[17][25] = 4'hD;
    SS8[18][25] = 4'hA;
    SS8[19][25] = 4'hA;
    SS8[20][25] = 4'hA;
    SS8[21][25] = 4'hD;
    SS8[22][25] = 4'hD;
    SS8[23][25] = 4'hD;
    SS8[24][25] = 4'hD;
    SS8[25][25] = 4'hC;
    SS8[26][25] = 4'hC;
    SS8[27][25] = 4'hC;
    SS8[28][25] = 4'hC;
    SS8[29][25] = 4'hC;
    SS8[30][25] = 4'hC;
    SS8[31][25] = 4'hC;
    SS8[32][25] = 4'hC;
    SS8[33][25] = 4'hC;
    SS8[34][25] = 4'hC;
    SS8[35][25] = 4'hC;
    SS8[36][25] = 4'hC;
    SS8[37][25] = 4'hC;
    SS8[38][25] = 4'hC;
    SS8[39][25] = 4'hD;
    SS8[40][25] = 4'h0;
    SS8[41][25] = 4'h0;
    SS8[42][25] = 4'h0;
    SS8[43][25] = 4'h0;
    SS8[44][25] = 4'h0;
    SS8[45][25] = 4'h0;
    SS8[46][25] = 4'h0;
    SS8[47][25] = 4'h0;
    SS8[0][26] = 4'h0;
    SS8[1][26] = 4'h0;
    SS8[2][26] = 4'h0;
    SS8[3][26] = 4'h0;
    SS8[4][26] = 4'h0;
    SS8[5][26] = 4'h0;
    SS8[6][26] = 4'h0;
    SS8[7][26] = 4'h0;
    SS8[8][26] = 4'h0;
    SS8[9][26] = 4'h0;
    SS8[10][26] = 4'h0;
    SS8[11][26] = 4'h0;
    SS8[12][26] = 4'h0;
    SS8[13][26] = 4'hD;
    SS8[14][26] = 4'hC;
    SS8[15][26] = 4'hC;
    SS8[16][26] = 4'hC;
    SS8[17][26] = 4'hC;
    SS8[18][26] = 4'hA;
    SS8[19][26] = 4'hA;
    SS8[20][26] = 4'hA;
    SS8[21][26] = 4'hA;
    SS8[22][26] = 4'hD;
    SS8[23][26] = 4'hD;
    SS8[24][26] = 4'hD;
    SS8[25][26] = 4'hD;
    SS8[26][26] = 4'hC;
    SS8[27][26] = 4'hC;
    SS8[28][26] = 4'hC;
    SS8[29][26] = 4'hC;
    SS8[30][26] = 4'hE;
    SS8[31][26] = 4'hC;
    SS8[32][26] = 4'hC;
    SS8[33][26] = 4'hC;
    SS8[34][26] = 4'hE;
    SS8[35][26] = 4'hC;
    SS8[36][26] = 4'hC;
    SS8[37][26] = 4'hC;
    SS8[38][26] = 4'hE;
    SS8[39][26] = 4'h0;
    SS8[40][26] = 4'h0;
    SS8[41][26] = 4'h0;
    SS8[42][26] = 4'h0;
    SS8[43][26] = 4'h0;
    SS8[44][26] = 4'h0;
    SS8[45][26] = 4'h0;
    SS8[46][26] = 4'h0;
    SS8[47][26] = 4'h0;
    SS8[0][27] = 4'h0;
    SS8[1][27] = 4'h0;
    SS8[2][27] = 4'h0;
    SS8[3][27] = 4'h0;
    SS8[4][27] = 4'h0;
    SS8[5][27] = 4'h0;
    SS8[6][27] = 4'h0;
    SS8[7][27] = 4'h0;
    SS8[8][27] = 4'h0;
    SS8[9][27] = 4'h0;
    SS8[10][27] = 4'h0;
    SS8[11][27] = 4'h0;
    SS8[12][27] = 4'hD;
    SS8[13][27] = 4'hD;
    SS8[14][27] = 4'hD;
    SS8[15][27] = 4'hC;
    SS8[16][27] = 4'hC;
    SS8[17][27] = 4'hC;
    SS8[18][27] = 4'hC;
    SS8[19][27] = 4'hA;
    SS8[20][27] = 4'hA;
    SS8[21][27] = 4'hA;
    SS8[22][27] = 4'hA;
    SS8[23][27] = 4'hD;
    SS8[24][27] = 4'hD;
    SS8[25][27] = 4'hC;
    SS8[26][27] = 4'hC;
    SS8[27][27] = 4'hC;
    SS8[28][27] = 4'hC;
    SS8[29][27] = 4'hE;
    SS8[30][27] = 4'hE;
    SS8[31][27] = 4'hE;
    SS8[32][27] = 4'hC;
    SS8[33][27] = 4'hE;
    SS8[34][27] = 4'hE;
    SS8[35][27] = 4'hE;
    SS8[36][27] = 4'hC;
    SS8[37][27] = 4'hE;
    SS8[38][27] = 4'hE;
    SS8[39][27] = 4'hE;
    SS8[40][27] = 4'h0;
    SS8[41][27] = 4'h0;
    SS8[42][27] = 4'h0;
    SS8[43][27] = 4'h0;
    SS8[44][27] = 4'h0;
    SS8[45][27] = 4'h0;
    SS8[46][27] = 4'h0;
    SS8[47][27] = 4'h0;
    SS8[0][28] = 4'h0;
    SS8[1][28] = 4'h0;
    SS8[2][28] = 4'h0;
    SS8[3][28] = 4'h0;
    SS8[4][28] = 4'h0;
    SS8[5][28] = 4'h0;
    SS8[6][28] = 4'h0;
    SS8[7][28] = 4'h0;
    SS8[8][28] = 4'h0;
    SS8[9][28] = 4'h0;
    SS8[10][28] = 4'h0;
    SS8[11][28] = 4'hD;
    SS8[12][28] = 4'hD;
    SS8[13][28] = 4'hD;
    SS8[14][28] = 4'hD;
    SS8[15][28] = 4'hC;
    SS8[16][28] = 4'hC;
    SS8[17][28] = 4'hC;
    SS8[18][28] = 4'hC;
    SS8[19][28] = 4'hC;
    SS8[20][28] = 4'hA;
    SS8[21][28] = 4'hA;
    SS8[22][28] = 4'hA;
    SS8[23][28] = 4'hA;
    SS8[24][28] = 4'hC;
    SS8[25][28] = 4'hC;
    SS8[26][28] = 4'hC;
    SS8[27][28] = 4'hC;
    SS8[28][28] = 4'hD;
    SS8[29][28] = 4'hE;
    SS8[30][28] = 4'hE;
    SS8[31][28] = 4'hE;
    SS8[32][28] = 4'hD;
    SS8[33][28] = 4'hE;
    SS8[34][28] = 4'hE;
    SS8[35][28] = 4'hE;
    SS8[36][28] = 4'hE;
    SS8[37][28] = 4'hE;
    SS8[38][28] = 4'hE;
    SS8[39][28] = 4'hE;
    SS8[40][28] = 4'hE;
    SS8[41][28] = 4'h0;
    SS8[42][28] = 4'h0;
    SS8[43][28] = 4'h0;
    SS8[44][28] = 4'h0;
    SS8[45][28] = 4'h0;
    SS8[46][28] = 4'h0;
    SS8[47][28] = 4'h0;
    SS8[0][29] = 4'h0;
    SS8[1][29] = 4'h0;
    SS8[2][29] = 4'h0;
    SS8[3][29] = 4'h0;
    SS8[4][29] = 4'h0;
    SS8[5][29] = 4'h0;
    SS8[6][29] = 4'h0;
    SS8[7][29] = 4'h0;
    SS8[8][29] = 4'h0;
    SS8[9][29] = 4'h0;
    SS8[10][29] = 4'hD;
    SS8[11][29] = 4'hD;
    SS8[12][29] = 4'hD;
    SS8[13][29] = 4'hD;
    SS8[14][29] = 4'hC;
    SS8[15][29] = 4'hC;
    SS8[16][29] = 4'hC;
    SS8[17][29] = 4'hC;
    SS8[18][29] = 4'hC;
    SS8[19][29] = 4'hC;
    SS8[20][29] = 4'hC;
    SS8[21][29] = 4'hA;
    SS8[22][29] = 4'hA;
    SS8[23][29] = 4'hD;
    SS8[24][29] = 4'hD;
    SS8[25][29] = 4'hC;
    SS8[26][29] = 4'hC;
    SS8[27][29] = 4'hD;
    SS8[28][29] = 4'hD;
    SS8[29][29] = 4'hD;
    SS8[30][29] = 4'hE;
    SS8[31][29] = 4'hD;
    SS8[32][29] = 4'hD;
    SS8[33][29] = 4'hD;
    SS8[34][29] = 4'hE;
    SS8[35][29] = 4'hE;
    SS8[36][29] = 4'hE;
    SS8[37][29] = 4'hE;
    SS8[38][29] = 4'hE;
    SS8[39][29] = 4'hE;
    SS8[40][29] = 4'hE;
    SS8[41][29] = 4'hE;
    SS8[42][29] = 4'h0;
    SS8[43][29] = 4'h0;
    SS8[44][29] = 4'h0;
    SS8[45][29] = 4'h0;
    SS8[46][29] = 4'h0;
    SS8[47][29] = 4'h0;
    SS8[0][30] = 4'h0;
    SS8[1][30] = 4'h0;
    SS8[2][30] = 4'h0;
    SS8[3][30] = 4'h0;
    SS8[4][30] = 4'h0;
    SS8[5][30] = 4'h0;
    SS8[6][30] = 4'h0;
    SS8[7][30] = 4'h0;
    SS8[8][30] = 4'h0;
    SS8[9][30] = 4'hD;
    SS8[10][30] = 4'hD;
    SS8[11][30] = 4'hD;
    SS8[12][30] = 4'hD;
    SS8[13][30] = 4'hC;
    SS8[14][30] = 4'hC;
    SS8[15][30] = 4'hC;
    SS8[16][30] = 4'hC;
    SS8[17][30] = 4'hC;
    SS8[18][30] = 4'hC;
    SS8[19][30] = 4'hC;
    SS8[20][30] = 4'hC;
    SS8[21][30] = 4'hC;
    SS8[22][30] = 4'hD;
    SS8[23][30] = 4'hD;
    SS8[24][30] = 4'hD;
    SS8[25][30] = 4'hD;
    SS8[26][30] = 4'hD;
    SS8[27][30] = 4'hD;
    SS8[28][30] = 4'hD;
    SS8[29][30] = 4'hD;
    SS8[30][30] = 4'hD;
    SS8[31][30] = 4'hD;
    SS8[32][30] = 4'hD;
    SS8[33][30] = 4'hD;
    SS8[34][30] = 4'hD;
    SS8[35][30] = 4'hE;
    SS8[36][30] = 4'hE;
    SS8[37][30] = 4'hE;
    SS8[38][30] = 4'hE;
    SS8[39][30] = 4'hE;
    SS8[40][30] = 4'hE;
    SS8[41][30] = 4'hE;
    SS8[42][30] = 4'hE;
    SS8[43][30] = 4'h0;
    SS8[44][30] = 4'h0;
    SS8[45][30] = 4'h0;
    SS8[46][30] = 4'h0;
    SS8[47][30] = 4'h0;
    SS8[0][31] = 4'h0;
    SS8[1][31] = 4'h0;
    SS8[2][31] = 4'h0;
    SS8[3][31] = 4'h0;
    SS8[4][31] = 4'h0;
    SS8[5][31] = 4'h0;
    SS8[6][31] = 4'h0;
    SS8[7][31] = 4'h0;
    SS8[8][31] = 4'hD;
    SS8[9][31] = 4'hD;
    SS8[10][31] = 4'hD;
    SS8[11][31] = 4'hD;
    SS8[12][31] = 4'hC;
    SS8[13][31] = 4'hC;
    SS8[14][31] = 4'hC;
    SS8[15][31] = 4'hC;
    SS8[16][31] = 4'hC;
    SS8[17][31] = 4'hC;
    SS8[18][31] = 4'hC;
    SS8[19][31] = 4'hC;
    SS8[20][31] = 4'hC;
    SS8[21][31] = 4'hC;
    SS8[22][31] = 4'hC;
    SS8[23][31] = 4'hD;
    SS8[24][31] = 4'hD;
    SS8[25][31] = 4'hD;
    SS8[26][31] = 4'hD;
    SS8[27][31] = 4'hD;
    SS8[28][31] = 4'hD;
    SS8[29][31] = 4'hD;
    SS8[30][31] = 4'hD;
    SS8[31][31] = 4'hD;
    SS8[32][31] = 4'hD;
    SS8[33][31] = 4'hD;
    SS8[34][31] = 4'hD;
    SS8[35][31] = 4'hD;
    SS8[36][31] = 4'hE;
    SS8[37][31] = 4'hE;
    SS8[38][31] = 4'hD;
    SS8[39][31] = 4'hD;
    SS8[40][31] = 4'hE;
    SS8[41][31] = 4'hE;
    SS8[42][31] = 4'hD;
    SS8[43][31] = 4'hD;
    SS8[44][31] = 4'h0;
    SS8[45][31] = 4'h0;
    SS8[46][31] = 4'h0;
    SS8[47][31] = 4'h0;
    SS8[0][32] = 4'h0;
    SS8[1][32] = 4'h0;
    SS8[2][32] = 4'h0;
    SS8[3][32] = 4'h0;
    SS8[4][32] = 4'h0;
    SS8[5][32] = 4'h0;
    SS8[6][32] = 4'h0;
    SS8[7][32] = 4'hD;
    SS8[8][32] = 4'hD;
    SS8[9][32] = 4'hD;
    SS8[10][32] = 4'hD;
    SS8[11][32] = 4'hC;
    SS8[12][32] = 4'hC;
    SS8[13][32] = 4'hC;
    SS8[14][32] = 4'hC;
    SS8[15][32] = 4'hC;
    SS8[16][32] = 4'hC;
    SS8[17][32] = 4'hC;
    SS8[18][32] = 4'hC;
    SS8[19][32] = 4'hC;
    SS8[20][32] = 4'hC;
    SS8[21][32] = 4'hC;
    SS8[22][32] = 4'hC;
    SS8[23][32] = 4'hC;
    SS8[24][32] = 4'hD;
    SS8[25][32] = 4'hD;
    SS8[26][32] = 4'hD;
    SS8[27][32] = 4'hD;
    SS8[28][32] = 4'hD;
    SS8[29][32] = 4'hD;
    SS8[30][32] = 4'hD;
    SS8[31][32] = 4'hD;
    SS8[32][32] = 4'hD;
    SS8[33][32] = 4'hD;
    SS8[34][32] = 4'hD;
    SS8[35][32] = 4'hD;
    SS8[36][32] = 4'hD;
    SS8[37][32] = 4'hD;
    SS8[38][32] = 4'hD;
    SS8[39][32] = 4'hD;
    SS8[40][32] = 4'hD;
    SS8[41][32] = 4'hD;
    SS8[42][32] = 4'hD;
    SS8[43][32] = 4'hD;
    SS8[44][32] = 4'hD;
    SS8[45][32] = 4'h0;
    SS8[46][32] = 4'h0;
    SS8[47][32] = 4'h0;
    SS8[0][33] = 4'h0;
    SS8[1][33] = 4'h0;
    SS8[2][33] = 4'h0;
    SS8[3][33] = 4'h0;
    SS8[4][33] = 4'h0;
    SS8[5][33] = 4'h0;
    SS8[6][33] = 4'h0;
    SS8[7][33] = 4'h0;
    SS8[8][33] = 4'hD;
    SS8[9][33] = 4'hD;
    SS8[10][33] = 4'hC;
    SS8[11][33] = 4'hC;
    SS8[12][33] = 4'hC;
    SS8[13][33] = 4'hC;
    SS8[14][33] = 4'hC;
    SS8[15][33] = 4'hC;
    SS8[16][33] = 4'hC;
    SS8[17][33] = 4'hC;
    SS8[18][33] = 4'hC;
    SS8[19][33] = 4'hD;
    SS8[20][33] = 4'hD;
    SS8[21][33] = 4'hC;
    SS8[22][33] = 4'hC;
    SS8[23][33] = 4'h0;
    SS8[24][33] = 4'h0;
    SS8[25][33] = 4'hD;
    SS8[26][33] = 4'hD;
    SS8[27][33] = 4'h3;
    SS8[28][33] = 4'h3;
    SS8[29][33] = 4'hD;
    SS8[30][33] = 4'hD;
    SS8[31][33] = 4'h0;
    SS8[32][33] = 4'h0;
    SS8[33][33] = 4'hE;
    SS8[34][33] = 4'hD;
    SS8[35][33] = 4'hD;
    SS8[36][33] = 4'h3;
    SS8[37][33] = 4'h3;
    SS8[38][33] = 4'hD;
    SS8[39][33] = 4'hD;
    SS8[40][33] = 4'hD;
    SS8[41][33] = 4'hD;
    SS8[42][33] = 4'hD;
    SS8[43][33] = 4'hD;
    SS8[44][33] = 4'hD;
    SS8[45][33] = 4'hD;
    SS8[46][33] = 4'h0;
    SS8[47][33] = 4'h0;
    SS8[0][34] = 4'h0;
    SS8[1][34] = 4'h0;
    SS8[2][34] = 4'h0;
    SS8[3][34] = 4'h0;
    SS8[4][34] = 4'h0;
    SS8[5][34] = 4'h0;
    SS8[6][34] = 4'h0;
    SS8[7][34] = 4'h0;
    SS8[8][34] = 4'h0;
    SS8[9][34] = 4'hC;
    SS8[10][34] = 4'hC;
    SS8[11][34] = 4'hC;
    SS8[12][34] = 4'hC;
    SS8[13][34] = 4'hC;
    SS8[14][34] = 4'hC;
    SS8[15][34] = 4'hC;
    SS8[16][34] = 4'hC;
    SS8[17][34] = 4'hC;
    SS8[18][34] = 4'hD;
    SS8[19][34] = 4'hD;
    SS8[20][34] = 4'hD;
    SS8[21][34] = 4'hD;
    SS8[22][34] = 4'h0;
    SS8[23][34] = 4'h0;
    SS8[24][34] = 4'h0;
    SS8[25][34] = 4'h0;
    SS8[26][34] = 4'h3;
    SS8[27][34] = 4'h3;
    SS8[28][34] = 4'h3;
    SS8[29][34] = 4'h3;
    SS8[30][34] = 4'h0;
    SS8[31][34] = 4'h0;
    SS8[32][34] = 4'h0;
    SS8[33][34] = 4'h0;
    SS8[34][34] = 4'hE;
    SS8[35][34] = 4'h3;
    SS8[36][34] = 4'h3;
    SS8[37][34] = 4'h3;
    SS8[38][34] = 4'h3;
    SS8[39][34] = 4'hD;
    SS8[40][34] = 4'hD;
    SS8[41][34] = 4'hD;
    SS8[42][34] = 4'hD;
    SS8[43][34] = 4'hD;
    SS8[44][34] = 4'hD;
    SS8[45][34] = 4'hD;
    SS8[46][34] = 4'hD;
    SS8[47][34] = 4'h0;
    SS8[0][35] = 4'h0;
    SS8[1][35] = 4'h0;
    SS8[2][35] = 4'h0;
    SS8[3][35] = 4'h0;
    SS8[4][35] = 4'h0;
    SS8[5][35] = 4'h0;
    SS8[6][35] = 4'h0;
    SS8[7][35] = 4'h0;
    SS8[8][35] = 4'hC;
    SS8[9][35] = 4'hC;
    SS8[10][35] = 4'hC;
    SS8[11][35] = 4'hC;
    SS8[12][35] = 4'hC;
    SS8[13][35] = 4'hC;
    SS8[14][35] = 4'hC;
    SS8[15][35] = 4'hC;
    SS8[16][35] = 4'hC;
    SS8[17][35] = 4'hD;
    SS8[18][35] = 4'hD;
    SS8[19][35] = 4'hD;
    SS8[20][35] = 4'hD;
    SS8[21][35] = 4'h0;
    SS8[22][35] = 4'h0;
    SS8[23][35] = 4'h0;
    SS8[24][35] = 4'h0;
    SS8[25][35] = 4'h0;
    SS8[26][35] = 4'h0;
    SS8[27][35] = 4'h3;
    SS8[28][35] = 4'h3;
    SS8[29][35] = 4'h2;
    SS8[30][35] = 4'h0;
    SS8[31][35] = 4'h0;
    SS8[32][35] = 4'h0;
    SS8[33][35] = 4'h0;
    SS8[34][35] = 4'h0;
    SS8[35][35] = 4'h2;
    SS8[36][35] = 4'h3;
    SS8[37][35] = 4'h3;
    SS8[38][35] = 4'h0;
    SS8[39][35] = 4'h0;
    SS8[40][35] = 4'hD;
    SS8[41][35] = 4'hD;
    SS8[42][35] = 4'h0;
    SS8[43][35] = 4'h0;
    SS8[44][35] = 4'hD;
    SS8[45][35] = 4'hD;
    SS8[46][35] = 4'h0;
    SS8[47][35] = 4'h0;
    SS8[0][36] = 4'h0;
    SS8[1][36] = 4'h0;
    SS8[2][36] = 4'h0;
    SS8[3][36] = 4'h0;
    SS8[4][36] = 4'h0;
    SS8[5][36] = 4'h0;
    SS8[6][36] = 4'h0;
    SS8[7][36] = 4'hC;
    SS8[8][36] = 4'hC;
    SS8[9][36] = 4'hC;
    SS8[10][36] = 4'hC;
    SS8[11][36] = 4'hC;
    SS8[12][36] = 4'hC;
    SS8[13][36] = 4'hC;
    SS8[14][36] = 4'hC;
    SS8[15][36] = 4'hC;
    SS8[16][36] = 4'hD;
    SS8[17][36] = 4'hD;
    SS8[18][36] = 4'hD;
    SS8[19][36] = 4'hD;
    SS8[20][36] = 4'h0;
    SS8[21][36] = 4'h0;
    SS8[22][36] = 4'h0;
    SS8[23][36] = 4'h0;
    SS8[24][36] = 4'h0;
    SS8[25][36] = 4'h0;
    SS8[26][36] = 4'h0;
    SS8[27][36] = 4'h0;
    SS8[28][36] = 4'h2;
    SS8[29][36] = 4'h0;
    SS8[30][36] = 4'h0;
    SS8[31][36] = 4'h0;
    SS8[32][36] = 4'h0;
    SS8[33][36] = 4'h0;
    SS8[34][36] = 4'h0;
    SS8[35][36] = 4'h0;
    SS8[36][36] = 4'h2;
    SS8[37][36] = 4'h0;
    SS8[38][36] = 4'h0;
    SS8[39][36] = 4'h0;
    SS8[40][36] = 4'h0;
    SS8[41][36] = 4'h0;
    SS8[42][36] = 4'h0;
    SS8[43][36] = 4'h0;
    SS8[44][36] = 4'h0;
    SS8[45][36] = 4'h0;
    SS8[46][36] = 4'h0;
    SS8[47][36] = 4'h0;
    SS8[0][37] = 4'h0;
    SS8[1][37] = 4'h0;
    SS8[2][37] = 4'h0;
    SS8[3][37] = 4'h0;
    SS8[4][37] = 4'h0;
    SS8[5][37] = 4'h0;
    SS8[6][37] = 4'hC;
    SS8[7][37] = 4'hC;
    SS8[8][37] = 4'hC;
    SS8[9][37] = 4'hC;
    SS8[10][37] = 4'hC;
    SS8[11][37] = 4'hC;
    SS8[12][37] = 4'hC;
    SS8[13][37] = 4'hC;
    SS8[14][37] = 4'hC;
    SS8[15][37] = 4'hD;
    SS8[16][37] = 4'hD;
    SS8[17][37] = 4'hD;
    SS8[18][37] = 4'hD;
    SS8[19][37] = 4'h0;
    SS8[20][37] = 4'h0;
    SS8[21][37] = 4'h0;
    SS8[22][37] = 4'h0;
    SS8[23][37] = 4'h0;
    SS8[24][37] = 4'h0;
    SS8[25][37] = 4'h0;
    SS8[26][37] = 4'h0;
    SS8[27][37] = 4'h0;
    SS8[28][37] = 4'h0;
    SS8[29][37] = 4'h0;
    SS8[30][37] = 4'h0;
    SS8[31][37] = 4'h0;
    SS8[32][37] = 4'h0;
    SS8[33][37] = 4'h0;
    SS8[34][37] = 4'h0;
    SS8[35][37] = 4'h0;
    SS8[36][37] = 4'h0;
    SS8[37][37] = 4'h0;
    SS8[38][37] = 4'h0;
    SS8[39][37] = 4'h0;
    SS8[40][37] = 4'h0;
    SS8[41][37] = 4'h0;
    SS8[42][37] = 4'h0;
    SS8[43][37] = 4'h0;
    SS8[44][37] = 4'h0;
    SS8[45][37] = 4'h0;
    SS8[46][37] = 4'h0;
    SS8[47][37] = 4'h0;
    SS8[0][38] = 4'h0;
    SS8[1][38] = 4'h0;
    SS8[2][38] = 4'h0;
    SS8[3][38] = 4'h0;
    SS8[4][38] = 4'h0;
    SS8[5][38] = 4'hC;
    SS8[6][38] = 4'hC;
    SS8[7][38] = 4'hC;
    SS8[8][38] = 4'hC;
    SS8[9][38] = 4'hC;
    SS8[10][38] = 4'hC;
    SS8[11][38] = 4'hC;
    SS8[12][38] = 4'hC;
    SS8[13][38] = 4'hC;
    SS8[14][38] = 4'hD;
    SS8[15][38] = 4'hD;
    SS8[16][38] = 4'hD;
    SS8[17][38] = 4'hD;
    SS8[18][38] = 4'h0;
    SS8[19][38] = 4'h0;
    SS8[20][38] = 4'h0;
    SS8[21][38] = 4'h0;
    SS8[22][38] = 4'h0;
    SS8[23][38] = 4'h0;
    SS8[24][38] = 4'h0;
    SS8[25][38] = 4'h0;
    SS8[26][38] = 4'h0;
    SS8[27][38] = 4'h0;
    SS8[28][38] = 4'h0;
    SS8[29][38] = 4'h0;
    SS8[30][38] = 4'h0;
    SS8[31][38] = 4'h0;
    SS8[32][38] = 4'h0;
    SS8[33][38] = 4'h0;
    SS8[34][38] = 4'h0;
    SS8[35][38] = 4'h0;
    SS8[36][38] = 4'h0;
    SS8[37][38] = 4'h0;
    SS8[38][38] = 4'h0;
    SS8[39][38] = 4'h0;
    SS8[40][38] = 4'h0;
    SS8[41][38] = 4'h0;
    SS8[42][38] = 4'h0;
    SS8[43][38] = 4'h0;
    SS8[44][38] = 4'h0;
    SS8[45][38] = 4'h0;
    SS8[46][38] = 4'h0;
    SS8[47][38] = 4'h0;
    SS8[0][39] = 4'h0;
    SS8[1][39] = 4'h0;
    SS8[2][39] = 4'h0;
    SS8[3][39] = 4'h0;
    SS8[4][39] = 4'h0;
    SS8[5][39] = 4'h0;
    SS8[6][39] = 4'hC;
    SS8[7][39] = 4'hC;
    SS8[8][39] = 4'hC;
    SS8[9][39] = 4'hC;
    SS8[10][39] = 4'hC;
    SS8[11][39] = 4'hC;
    SS8[12][39] = 4'hC;
    SS8[13][39] = 4'h0;
    SS8[14][39] = 4'hD;
    SS8[15][39] = 4'hD;
    SS8[16][39] = 4'hD;
    SS8[17][39] = 4'h0;
    SS8[18][39] = 4'h0;
    SS8[19][39] = 4'h0;
    SS8[20][39] = 4'h0;
    SS8[21][39] = 4'h0;
    SS8[22][39] = 4'h0;
    SS8[23][39] = 4'h0;
    SS8[24][39] = 4'h0;
    SS8[25][39] = 4'h0;
    SS8[26][39] = 4'h0;
    SS8[27][39] = 4'h0;
    SS8[28][39] = 4'h0;
    SS8[29][39] = 4'h0;
    SS8[30][39] = 4'h0;
    SS8[31][39] = 4'h0;
    SS8[32][39] = 4'h0;
    SS8[33][39] = 4'h0;
    SS8[34][39] = 4'h0;
    SS8[35][39] = 4'h0;
    SS8[36][39] = 4'h0;
    SS8[37][39] = 4'h0;
    SS8[38][39] = 4'h0;
    SS8[39][39] = 4'h0;
    SS8[40][39] = 4'h0;
    SS8[41][39] = 4'h0;
    SS8[42][39] = 4'h0;
    SS8[43][39] = 4'h0;
    SS8[44][39] = 4'h0;
    SS8[45][39] = 4'h0;
    SS8[46][39] = 4'h0;
    SS8[47][39] = 4'h0;
    SS8[0][40] = 4'h0;
    SS8[1][40] = 4'h0;
    SS8[2][40] = 4'h0;
    SS8[3][40] = 4'h0;
    SS8[4][40] = 4'h0;
    SS8[5][40] = 4'h0;
    SS8[6][40] = 4'h0;
    SS8[7][40] = 4'hC;
    SS8[8][40] = 4'hC;
    SS8[9][40] = 4'hC;
    SS8[10][40] = 4'hC;
    SS8[11][40] = 4'hC;
    SS8[12][40] = 4'h0;
    SS8[13][40] = 4'h0;
    SS8[14][40] = 4'h0;
    SS8[15][40] = 4'hD;
    SS8[16][40] = 4'h0;
    SS8[17][40] = 4'h0;
    SS8[18][40] = 4'h0;
    SS8[19][40] = 4'h0;
    SS8[20][40] = 4'h0;
    SS8[21][40] = 4'h0;
    SS8[22][40] = 4'h0;
    SS8[23][40] = 4'h0;
    SS8[24][40] = 4'h0;
    SS8[25][40] = 4'h0;
    SS8[26][40] = 4'h0;
    SS8[27][40] = 4'h0;
    SS8[28][40] = 4'h0;
    SS8[29][40] = 4'h0;
    SS8[30][40] = 4'h0;
    SS8[31][40] = 4'h0;
    SS8[32][40] = 4'h0;
    SS8[33][40] = 4'h0;
    SS8[34][40] = 4'h0;
    SS8[35][40] = 4'h0;
    SS8[36][40] = 4'h0;
    SS8[37][40] = 4'h0;
    SS8[38][40] = 4'h0;
    SS8[39][40] = 4'h0;
    SS8[40][40] = 4'h0;
    SS8[41][40] = 4'h0;
    SS8[42][40] = 4'h0;
    SS8[43][40] = 4'h0;
    SS8[44][40] = 4'h0;
    SS8[45][40] = 4'h0;
    SS8[46][40] = 4'h0;
    SS8[47][40] = 4'h0;
    SS8[0][41] = 4'h0;
    SS8[1][41] = 4'h0;
    SS8[2][41] = 4'h0;
    SS8[3][41] = 4'h0;
    SS8[4][41] = 4'h0;
    SS8[5][41] = 4'h0;
    SS8[6][41] = 4'h0;
    SS8[7][41] = 4'h0;
    SS8[8][41] = 4'hC;
    SS8[9][41] = 4'hC;
    SS8[10][41] = 4'hC;
    SS8[11][41] = 4'h0;
    SS8[12][41] = 4'h0;
    SS8[13][41] = 4'h0;
    SS8[14][41] = 4'h0;
    SS8[15][41] = 4'h0;
    SS8[16][41] = 4'h0;
    SS8[17][41] = 4'h0;
    SS8[18][41] = 4'h0;
    SS8[19][41] = 4'h0;
    SS8[20][41] = 4'h0;
    SS8[21][41] = 4'h0;
    SS8[22][41] = 4'h0;
    SS8[23][41] = 4'h0;
    SS8[24][41] = 4'h0;
    SS8[25][41] = 4'h0;
    SS8[26][41] = 4'h0;
    SS8[27][41] = 4'h0;
    SS8[28][41] = 4'h0;
    SS8[29][41] = 4'h0;
    SS8[30][41] = 4'h0;
    SS8[31][41] = 4'h0;
    SS8[32][41] = 4'h0;
    SS8[33][41] = 4'h0;
    SS8[34][41] = 4'h0;
    SS8[35][41] = 4'h0;
    SS8[36][41] = 4'h0;
    SS8[37][41] = 4'h0;
    SS8[38][41] = 4'h0;
    SS8[39][41] = 4'h0;
    SS8[40][41] = 4'h0;
    SS8[41][41] = 4'h0;
    SS8[42][41] = 4'h0;
    SS8[43][41] = 4'h0;
    SS8[44][41] = 4'h0;
    SS8[45][41] = 4'h0;
    SS8[46][41] = 4'h0;
    SS8[47][41] = 4'h0;
    SS8[0][42] = 4'h0;
    SS8[1][42] = 4'h0;
    SS8[2][42] = 4'h0;
    SS8[3][42] = 4'h0;
    SS8[4][42] = 4'h0;
    SS8[5][42] = 4'h0;
    SS8[6][42] = 4'h0;
    SS8[7][42] = 4'h0;
    SS8[8][42] = 4'h0;
    SS8[9][42] = 4'hC;
    SS8[10][42] = 4'h0;
    SS8[11][42] = 4'h0;
    SS8[12][42] = 4'h0;
    SS8[13][42] = 4'h0;
    SS8[14][42] = 4'h0;
    SS8[15][42] = 4'h0;
    SS8[16][42] = 4'h0;
    SS8[17][42] = 4'h0;
    SS8[18][42] = 4'h0;
    SS8[19][42] = 4'h0;
    SS8[20][42] = 4'h0;
    SS8[21][42] = 4'h0;
    SS8[22][42] = 4'h0;
    SS8[23][42] = 4'h0;
    SS8[24][42] = 4'h0;
    SS8[25][42] = 4'h0;
    SS8[26][42] = 4'h0;
    SS8[27][42] = 4'h0;
    SS8[28][42] = 4'h0;
    SS8[29][42] = 4'h0;
    SS8[30][42] = 4'h0;
    SS8[31][42] = 4'h0;
    SS8[32][42] = 4'h0;
    SS8[33][42] = 4'h0;
    SS8[34][42] = 4'h0;
    SS8[35][42] = 4'h0;
    SS8[36][42] = 4'h0;
    SS8[37][42] = 4'h0;
    SS8[38][42] = 4'h0;
    SS8[39][42] = 4'h0;
    SS8[40][42] = 4'h0;
    SS8[41][42] = 4'h0;
    SS8[42][42] = 4'h0;
    SS8[43][42] = 4'h0;
    SS8[44][42] = 4'h0;
    SS8[45][42] = 4'h0;
    SS8[46][42] = 4'h0;
    SS8[47][42] = 4'h0;
    SS8[0][43] = 4'h0;
    SS8[1][43] = 4'h0;
    SS8[2][43] = 4'h0;
    SS8[3][43] = 4'h0;
    SS8[4][43] = 4'h0;
    SS8[5][43] = 4'h0;
    SS8[6][43] = 4'h0;
    SS8[7][43] = 4'h0;
    SS8[8][43] = 4'h0;
    SS8[9][43] = 4'h0;
    SS8[10][43] = 4'h0;
    SS8[11][43] = 4'h0;
    SS8[12][43] = 4'h0;
    SS8[13][43] = 4'h0;
    SS8[14][43] = 4'h0;
    SS8[15][43] = 4'h0;
    SS8[16][43] = 4'h0;
    SS8[17][43] = 4'h0;
    SS8[18][43] = 4'h0;
    SS8[19][43] = 4'h0;
    SS8[20][43] = 4'h0;
    SS8[21][43] = 4'h0;
    SS8[22][43] = 4'h0;
    SS8[23][43] = 4'h0;
    SS8[24][43] = 4'h0;
    SS8[25][43] = 4'h0;
    SS8[26][43] = 4'h0;
    SS8[27][43] = 4'h0;
    SS8[28][43] = 4'h0;
    SS8[29][43] = 4'h0;
    SS8[30][43] = 4'h0;
    SS8[31][43] = 4'h0;
    SS8[32][43] = 4'h0;
    SS8[33][43] = 4'h0;
    SS8[34][43] = 4'h0;
    SS8[35][43] = 4'h0;
    SS8[36][43] = 4'h0;
    SS8[37][43] = 4'h0;
    SS8[38][43] = 4'h0;
    SS8[39][43] = 4'h0;
    SS8[40][43] = 4'h0;
    SS8[41][43] = 4'h0;
    SS8[42][43] = 4'h0;
    SS8[43][43] = 4'h0;
    SS8[44][43] = 4'h0;
    SS8[45][43] = 4'h0;
    SS8[46][43] = 4'h0;
    SS8[47][43] = 4'h0;
    SS8[0][44] = 4'h0;
    SS8[1][44] = 4'h0;
    SS8[2][44] = 4'h0;
    SS8[3][44] = 4'h0;
    SS8[4][44] = 4'h0;
    SS8[5][44] = 4'h0;
    SS8[6][44] = 4'h0;
    SS8[7][44] = 4'h0;
    SS8[8][44] = 4'h0;
    SS8[9][44] = 4'h0;
    SS8[10][44] = 4'h0;
    SS8[11][44] = 4'h0;
    SS8[12][44] = 4'h0;
    SS8[13][44] = 4'h0;
    SS8[14][44] = 4'h0;
    SS8[15][44] = 4'h0;
    SS8[16][44] = 4'h0;
    SS8[17][44] = 4'h0;
    SS8[18][44] = 4'h0;
    SS8[19][44] = 4'h0;
    SS8[20][44] = 4'h0;
    SS8[21][44] = 4'h0;
    SS8[22][44] = 4'h0;
    SS8[23][44] = 4'h0;
    SS8[24][44] = 4'h0;
    SS8[25][44] = 4'h0;
    SS8[26][44] = 4'h0;
    SS8[27][44] = 4'h0;
    SS8[28][44] = 4'h0;
    SS8[29][44] = 4'h0;
    SS8[30][44] = 4'h0;
    SS8[31][44] = 4'h0;
    SS8[32][44] = 4'h0;
    SS8[33][44] = 4'h0;
    SS8[34][44] = 4'h0;
    SS8[35][44] = 4'h0;
    SS8[36][44] = 4'h0;
    SS8[37][44] = 4'h0;
    SS8[38][44] = 4'h0;
    SS8[39][44] = 4'h0;
    SS8[40][44] = 4'h0;
    SS8[41][44] = 4'h0;
    SS8[42][44] = 4'h0;
    SS8[43][44] = 4'h0;
    SS8[44][44] = 4'h0;
    SS8[45][44] = 4'h0;
    SS8[46][44] = 4'h0;
    SS8[47][44] = 4'h0;
    SS8[0][45] = 4'h0;
    SS8[1][45] = 4'h0;
    SS8[2][45] = 4'h0;
    SS8[3][45] = 4'h0;
    SS8[4][45] = 4'h0;
    SS8[5][45] = 4'h0;
    SS8[6][45] = 4'h0;
    SS8[7][45] = 4'h0;
    SS8[8][45] = 4'h0;
    SS8[9][45] = 4'h0;
    SS8[10][45] = 4'h0;
    SS8[11][45] = 4'h0;
    SS8[12][45] = 4'h0;
    SS8[13][45] = 4'h0;
    SS8[14][45] = 4'h0;
    SS8[15][45] = 4'h0;
    SS8[16][45] = 4'h0;
    SS8[17][45] = 4'h0;
    SS8[18][45] = 4'h0;
    SS8[19][45] = 4'h0;
    SS8[20][45] = 4'h0;
    SS8[21][45] = 4'h0;
    SS8[22][45] = 4'h0;
    SS8[23][45] = 4'h0;
    SS8[24][45] = 4'h0;
    SS8[25][45] = 4'h0;
    SS8[26][45] = 4'h0;
    SS8[27][45] = 4'h0;
    SS8[28][45] = 4'h0;
    SS8[29][45] = 4'h0;
    SS8[30][45] = 4'h0;
    SS8[31][45] = 4'h0;
    SS8[32][45] = 4'h0;
    SS8[33][45] = 4'h0;
    SS8[34][45] = 4'h0;
    SS8[35][45] = 4'h0;
    SS8[36][45] = 4'h0;
    SS8[37][45] = 4'h0;
    SS8[38][45] = 4'h0;
    SS8[39][45] = 4'h0;
    SS8[40][45] = 4'h0;
    SS8[41][45] = 4'h0;
    SS8[42][45] = 4'h0;
    SS8[43][45] = 4'h0;
    SS8[44][45] = 4'h0;
    SS8[45][45] = 4'h0;
    SS8[46][45] = 4'h0;
    SS8[47][45] = 4'h0;
    SS8[0][46] = 4'h0;
    SS8[1][46] = 4'h0;
    SS8[2][46] = 4'h0;
    SS8[3][46] = 4'h0;
    SS8[4][46] = 4'h0;
    SS8[5][46] = 4'h0;
    SS8[6][46] = 4'h0;
    SS8[7][46] = 4'h0;
    SS8[8][46] = 4'h0;
    SS8[9][46] = 4'h0;
    SS8[10][46] = 4'h0;
    SS8[11][46] = 4'h0;
    SS8[12][46] = 4'h0;
    SS8[13][46] = 4'h0;
    SS8[14][46] = 4'h0;
    SS8[15][46] = 4'h0;
    SS8[16][46] = 4'h0;
    SS8[17][46] = 4'h0;
    SS8[18][46] = 4'h0;
    SS8[19][46] = 4'h0;
    SS8[20][46] = 4'h0;
    SS8[21][46] = 4'h0;
    SS8[22][46] = 4'h0;
    SS8[23][46] = 4'h0;
    SS8[24][46] = 4'h0;
    SS8[25][46] = 4'h0;
    SS8[26][46] = 4'h0;
    SS8[27][46] = 4'h0;
    SS8[28][46] = 4'h0;
    SS8[29][46] = 4'h0;
    SS8[30][46] = 4'h0;
    SS8[31][46] = 4'h0;
    SS8[32][46] = 4'h0;
    SS8[33][46] = 4'h0;
    SS8[34][46] = 4'h0;
    SS8[35][46] = 4'h0;
    SS8[36][46] = 4'h0;
    SS8[37][46] = 4'h0;
    SS8[38][46] = 4'h0;
    SS8[39][46] = 4'h0;
    SS8[40][46] = 4'h0;
    SS8[41][46] = 4'h0;
    SS8[42][46] = 4'h0;
    SS8[43][46] = 4'h0;
    SS8[44][46] = 4'h0;
    SS8[45][46] = 4'h0;
    SS8[46][46] = 4'h0;
    SS8[47][46] = 4'h0;
    SS8[0][47] = 4'h0;
    SS8[1][47] = 4'h0;
    SS8[2][47] = 4'h0;
    SS8[3][47] = 4'h0;
    SS8[4][47] = 4'h0;
    SS8[5][47] = 4'h0;
    SS8[6][47] = 4'h0;
    SS8[7][47] = 4'h0;
    SS8[8][47] = 4'h0;
    SS8[9][47] = 4'h0;
    SS8[10][47] = 4'h0;
    SS8[11][47] = 4'h0;
    SS8[12][47] = 4'h0;
    SS8[13][47] = 4'h0;
    SS8[14][47] = 4'h0;
    SS8[15][47] = 4'h0;
    SS8[16][47] = 4'h0;
    SS8[17][47] = 4'h0;
    SS8[18][47] = 4'h0;
    SS8[19][47] = 4'h0;
    SS8[20][47] = 4'h0;
    SS8[21][47] = 4'h0;
    SS8[22][47] = 4'h0;
    SS8[23][47] = 4'h0;
    SS8[24][47] = 4'h0;
    SS8[25][47] = 4'h0;
    SS8[26][47] = 4'h0;
    SS8[27][47] = 4'h0;
    SS8[28][47] = 4'h0;
    SS8[29][47] = 4'h0;
    SS8[30][47] = 4'h0;
    SS8[31][47] = 4'h0;
    SS8[32][47] = 4'h0;
    SS8[33][47] = 4'h0;
    SS8[34][47] = 4'h0;
    SS8[35][47] = 4'h0;
    SS8[36][47] = 4'h0;
    SS8[37][47] = 4'h0;
    SS8[38][47] = 4'h0;
    SS8[39][47] = 4'h0;
    SS8[40][47] = 4'h0;
    SS8[41][47] = 4'h0;
    SS8[42][47] = 4'h0;
    SS8[43][47] = 4'h0;
    SS8[44][47] = 4'h0;
    SS8[45][47] = 4'h0;
    SS8[46][47] = 4'h0;
    SS8[47][47] = 4'h0;
 
//SS 9
    SS9[0][0] = 4'h0;
    SS9[1][0] = 4'h0;
    SS9[2][0] = 4'h0;
    SS9[3][0] = 4'h0;
    SS9[4][0] = 4'h0;
    SS9[5][0] = 4'h0;
    SS9[6][0] = 4'h0;
    SS9[7][0] = 4'h0;
    SS9[8][0] = 4'h0;
    SS9[9][0] = 4'h0;
    SS9[10][0] = 4'h0;
    SS9[11][0] = 4'h0;
    SS9[12][0] = 4'h0;
    SS9[13][0] = 4'h0;
    SS9[14][0] = 4'h0;
    SS9[15][0] = 4'h0;
    SS9[16][0] = 4'h0;
    SS9[17][0] = 4'h0;
    SS9[18][0] = 4'h0;
    SS9[19][0] = 4'h0;
    SS9[20][0] = 4'h0;
    SS9[21][0] = 4'hD;
    SS9[22][0] = 4'hD;
    SS9[23][0] = 4'hD;
    SS9[24][0] = 4'h0;
    SS9[25][0] = 4'h0;
    SS9[26][0] = 4'h0;
    SS9[27][0] = 4'h0;
    SS9[28][0] = 4'h0;
    SS9[29][0] = 4'h0;
    SS9[30][0] = 4'h0;
    SS9[31][0] = 4'h0;
    SS9[32][0] = 4'h0;
    SS9[33][0] = 4'h0;
    SS9[34][0] = 4'h0;
    SS9[35][0] = 4'h0;
    SS9[36][0] = 4'h0;
    SS9[37][0] = 4'h0;
    SS9[38][0] = 4'h0;
    SS9[39][0] = 4'h0;
    SS9[40][0] = 4'h0;
    SS9[41][0] = 4'h0;
    SS9[42][0] = 4'h0;
    SS9[43][0] = 4'h0;
    SS9[44][0] = 4'h0;
    SS9[45][0] = 4'h0;
    SS9[46][0] = 4'h0;
    SS9[47][0] = 4'h0;
    SS9[0][1] = 4'h0;
    SS9[1][1] = 4'h0;
    SS9[2][1] = 4'h0;
    SS9[3][1] = 4'h0;
    SS9[4][1] = 4'h0;
    SS9[5][1] = 4'h0;
    SS9[6][1] = 4'h0;
    SS9[7][1] = 4'h0;
    SS9[8][1] = 4'h0;
    SS9[9][1] = 4'h0;
    SS9[10][1] = 4'h0;
    SS9[11][1] = 4'h0;
    SS9[12][1] = 4'h0;
    SS9[13][1] = 4'h0;
    SS9[14][1] = 4'h0;
    SS9[15][1] = 4'h0;
    SS9[16][1] = 4'h0;
    SS9[17][1] = 4'h0;
    SS9[18][1] = 4'h0;
    SS9[19][1] = 4'h0;
    SS9[20][1] = 4'h0;
    SS9[21][1] = 4'hD;
    SS9[22][1] = 4'hD;
    SS9[23][1] = 4'hD;
    SS9[24][1] = 4'h0;
    SS9[25][1] = 4'h0;
    SS9[26][1] = 4'h0;
    SS9[27][1] = 4'h0;
    SS9[28][1] = 4'h0;
    SS9[29][1] = 4'h0;
    SS9[30][1] = 4'h0;
    SS9[31][1] = 4'h0;
    SS9[32][1] = 4'h0;
    SS9[33][1] = 4'h0;
    SS9[34][1] = 4'h0;
    SS9[35][1] = 4'h0;
    SS9[36][1] = 4'h0;
    SS9[37][1] = 4'h0;
    SS9[38][1] = 4'h0;
    SS9[39][1] = 4'h0;
    SS9[40][1] = 4'h0;
    SS9[41][1] = 4'h0;
    SS9[42][1] = 4'h0;
    SS9[43][1] = 4'h0;
    SS9[44][1] = 4'h0;
    SS9[45][1] = 4'h0;
    SS9[46][1] = 4'h0;
    SS9[47][1] = 4'h0;
    SS9[0][2] = 4'h0;
    SS9[1][2] = 4'h0;
    SS9[2][2] = 4'h0;
    SS9[3][2] = 4'h0;
    SS9[4][2] = 4'h0;
    SS9[5][2] = 4'h0;
    SS9[6][2] = 4'h0;
    SS9[7][2] = 4'h0;
    SS9[8][2] = 4'h0;
    SS9[9][2] = 4'h0;
    SS9[10][2] = 4'h0;
    SS9[11][2] = 4'h0;
    SS9[12][2] = 4'h0;
    SS9[13][2] = 4'h0;
    SS9[14][2] = 4'h0;
    SS9[15][2] = 4'h0;
    SS9[16][2] = 4'h0;
    SS9[17][2] = 4'h0;
    SS9[18][2] = 4'h0;
    SS9[19][2] = 4'h0;
    SS9[20][2] = 4'h0;
    SS9[21][2] = 4'hE;
    SS9[22][2] = 4'hD;
    SS9[23][2] = 4'hD;
    SS9[24][2] = 4'hD;
    SS9[25][2] = 4'h0;
    SS9[26][2] = 4'h0;
    SS9[27][2] = 4'h0;
    SS9[28][2] = 4'h0;
    SS9[29][2] = 4'h0;
    SS9[30][2] = 4'h0;
    SS9[31][2] = 4'h0;
    SS9[32][2] = 4'h0;
    SS9[33][2] = 4'h0;
    SS9[34][2] = 4'h0;
    SS9[35][2] = 4'h0;
    SS9[36][2] = 4'h0;
    SS9[37][2] = 4'hC;
    SS9[38][2] = 4'hD;
    SS9[39][2] = 4'hD;
    SS9[40][2] = 4'hD;
    SS9[41][2] = 4'h0;
    SS9[42][2] = 4'h0;
    SS9[43][2] = 4'h0;
    SS9[44][2] = 4'h0;
    SS9[45][2] = 4'h0;
    SS9[46][2] = 4'h0;
    SS9[47][2] = 4'h0;
    SS9[0][3] = 4'h0;
    SS9[1][3] = 4'h0;
    SS9[2][3] = 4'h0;
    SS9[3][3] = 4'h0;
    SS9[4][3] = 4'h0;
    SS9[5][3] = 4'h0;
    SS9[6][3] = 4'h0;
    SS9[7][3] = 4'h0;
    SS9[8][3] = 4'h0;
    SS9[9][3] = 4'h0;
    SS9[10][3] = 4'h0;
    SS9[11][3] = 4'h0;
    SS9[12][3] = 4'h0;
    SS9[13][3] = 4'h0;
    SS9[14][3] = 4'h0;
    SS9[15][3] = 4'h0;
    SS9[16][3] = 4'h0;
    SS9[17][3] = 4'h0;
    SS9[18][3] = 4'h0;
    SS9[19][3] = 4'hD;
    SS9[20][3] = 4'hD;
    SS9[21][3] = 4'hD;
    SS9[22][3] = 4'hD;
    SS9[23][3] = 4'hD;
    SS9[24][3] = 4'hD;
    SS9[25][3] = 4'h0;
    SS9[26][3] = 4'h0;
    SS9[27][3] = 4'h0;
    SS9[28][3] = 4'h0;
    SS9[29][3] = 4'h0;
    SS9[30][3] = 4'h0;
    SS9[31][3] = 4'h0;
    SS9[32][3] = 4'h0;
    SS9[33][3] = 4'h0;
    SS9[34][3] = 4'h0;
    SS9[35][3] = 4'hC;
    SS9[36][3] = 4'hC;
    SS9[37][3] = 4'hC;
    SS9[38][3] = 4'hD;
    SS9[39][3] = 4'hD;
    SS9[40][3] = 4'hD;
    SS9[41][3] = 4'h0;
    SS9[42][3] = 4'h0;
    SS9[43][3] = 4'h0;
    SS9[44][3] = 4'h0;
    SS9[45][3] = 4'h0;
    SS9[46][3] = 4'h0;
    SS9[47][3] = 4'h0;
    SS9[0][4] = 4'h0;
    SS9[1][4] = 4'h0;
    SS9[2][4] = 4'h0;
    SS9[3][4] = 4'h0;
    SS9[4][4] = 4'h0;
    SS9[5][4] = 4'h0;
    SS9[6][4] = 4'h0;
    SS9[7][4] = 4'h0;
    SS9[8][4] = 4'h0;
    SS9[9][4] = 4'h0;
    SS9[10][4] = 4'h0;
    SS9[11][4] = 4'h0;
    SS9[12][4] = 4'h0;
    SS9[13][4] = 4'h0;
    SS9[14][4] = 4'h0;
    SS9[15][4] = 4'h0;
    SS9[16][4] = 4'h0;
    SS9[17][4] = 4'h0;
    SS9[18][4] = 4'h0;
    SS9[19][4] = 4'hD;
    SS9[20][4] = 4'hD;
    SS9[21][4] = 4'hD;
    SS9[22][4] = 4'hD;
    SS9[23][4] = 4'hD;
    SS9[24][4] = 4'hD;
    SS9[25][4] = 4'hE;
    SS9[26][4] = 4'h0;
    SS9[27][4] = 4'h0;
    SS9[28][4] = 4'h0;
    SS9[29][4] = 4'h0;
    SS9[30][4] = 4'h0;
    SS9[31][4] = 4'h0;
    SS9[32][4] = 4'hC;
    SS9[33][4] = 4'hC;
    SS9[34][4] = 4'hC;
    SS9[35][4] = 4'hC;
    SS9[36][4] = 4'hC;
    SS9[37][4] = 4'hC;
    SS9[38][4] = 4'hD;
    SS9[39][4] = 4'hD;
    SS9[40][4] = 4'h0;
    SS9[41][4] = 4'h0;
    SS9[42][4] = 4'h0;
    SS9[43][4] = 4'h0;
    SS9[44][4] = 4'h0;
    SS9[45][4] = 4'h0;
    SS9[46][4] = 4'h0;
    SS9[47][4] = 4'h0;
    SS9[0][5] = 4'h0;
    SS9[1][5] = 4'h0;
    SS9[2][5] = 4'h0;
    SS9[3][5] = 4'h0;
    SS9[4][5] = 4'h0;
    SS9[5][5] = 4'h0;
    SS9[6][5] = 4'h0;
    SS9[7][5] = 4'h0;
    SS9[8][5] = 4'h0;
    SS9[9][5] = 4'h0;
    SS9[10][5] = 4'h0;
    SS9[11][5] = 4'h0;
    SS9[12][5] = 4'h0;
    SS9[13][5] = 4'h0;
    SS9[14][5] = 4'h0;
    SS9[15][5] = 4'h0;
    SS9[16][5] = 4'h0;
    SS9[17][5] = 4'h0;
    SS9[18][5] = 4'h0;
    SS9[19][5] = 4'h0;
    SS9[20][5] = 4'hD;
    SS9[21][5] = 4'hD;
    SS9[22][5] = 4'hD;
    SS9[23][5] = 4'hE;
    SS9[24][5] = 4'hE;
    SS9[25][5] = 4'hE;
    SS9[26][5] = 4'h0;
    SS9[27][5] = 4'h0;
    SS9[28][5] = 4'h0;
    SS9[29][5] = 4'h0;
    SS9[30][5] = 4'h0;
    SS9[31][5] = 4'h0;
    SS9[32][5] = 4'hC;
    SS9[33][5] = 4'hC;
    SS9[34][5] = 4'hC;
    SS9[35][5] = 4'hC;
    SS9[36][5] = 4'hC;
    SS9[37][5] = 4'hC;
    SS9[38][5] = 4'hD;
    SS9[39][5] = 4'h0;
    SS9[40][5] = 4'h0;
    SS9[41][5] = 4'h0;
    SS9[42][5] = 4'h0;
    SS9[43][5] = 4'h0;
    SS9[44][5] = 4'h0;
    SS9[45][5] = 4'h0;
    SS9[46][5] = 4'h0;
    SS9[47][5] = 4'h0;
    SS9[0][6] = 4'h0;
    SS9[1][6] = 4'h0;
    SS9[2][6] = 4'h0;
    SS9[3][6] = 4'h0;
    SS9[4][6] = 4'h0;
    SS9[5][6] = 4'h0;
    SS9[6][6] = 4'h0;
    SS9[7][6] = 4'h0;
    SS9[8][6] = 4'h0;
    SS9[9][6] = 4'h0;
    SS9[10][6] = 4'h0;
    SS9[11][6] = 4'h0;
    SS9[12][6] = 4'h0;
    SS9[13][6] = 4'h0;
    SS9[14][6] = 4'h0;
    SS9[15][6] = 4'h0;
    SS9[16][6] = 4'h0;
    SS9[17][6] = 4'h0;
    SS9[18][6] = 4'h0;
    SS9[19][6] = 4'h0;
    SS9[20][6] = 4'hD;
    SS9[21][6] = 4'hD;
    SS9[22][6] = 4'hD;
    SS9[23][6] = 4'hE;
    SS9[24][6] = 4'hE;
    SS9[25][6] = 4'hE;
    SS9[26][6] = 4'h0;
    SS9[27][6] = 4'h0;
    SS9[28][6] = 4'h0;
    SS9[29][6] = 4'h0;
    SS9[30][6] = 4'h0;
    SS9[31][6] = 4'h0;
    SS9[32][6] = 4'h0;
    SS9[33][6] = 4'hC;
    SS9[34][6] = 4'hC;
    SS9[35][6] = 4'hC;
    SS9[36][6] = 4'hD;
    SS9[37][6] = 4'hD;
    SS9[38][6] = 4'hD;
    SS9[39][6] = 4'h0;
    SS9[40][6] = 4'h0;
    SS9[41][6] = 4'h0;
    SS9[42][6] = 4'h0;
    SS9[43][6] = 4'h0;
    SS9[44][6] = 4'h0;
    SS9[45][6] = 4'h0;
    SS9[46][6] = 4'h0;
    SS9[47][6] = 4'h0;
    SS9[0][7] = 4'h0;
    SS9[1][7] = 4'h0;
    SS9[2][7] = 4'h0;
    SS9[3][7] = 4'h0;
    SS9[4][7] = 4'h0;
    SS9[5][7] = 4'h0;
    SS9[6][7] = 4'h0;
    SS9[7][7] = 4'h0;
    SS9[8][7] = 4'h0;
    SS9[9][7] = 4'h0;
    SS9[10][7] = 4'h0;
    SS9[11][7] = 4'h0;
    SS9[12][7] = 4'h0;
    SS9[13][7] = 4'h0;
    SS9[14][7] = 4'h0;
    SS9[15][7] = 4'h0;
    SS9[16][7] = 4'h0;
    SS9[17][7] = 4'h3;
    SS9[18][7] = 4'h3;
    SS9[19][7] = 4'h3;
    SS9[20][7] = 4'hD;
    SS9[21][7] = 4'hD;
    SS9[22][7] = 4'hD;
    SS9[23][7] = 4'hD;
    SS9[24][7] = 4'hE;
    SS9[25][7] = 4'hE;
    SS9[26][7] = 4'hE;
    SS9[27][7] = 4'h0;
    SS9[28][7] = 4'h0;
    SS9[29][7] = 4'h0;
    SS9[30][7] = 4'h0;
    SS9[31][7] = 4'h0;
    SS9[32][7] = 4'h0;
    SS9[33][7] = 4'hC;
    SS9[34][7] = 4'hC;
    SS9[35][7] = 4'hC;
    SS9[36][7] = 4'hD;
    SS9[37][7] = 4'hD;
    SS9[38][7] = 4'hD;
    SS9[39][7] = 4'hD;
    SS9[40][7] = 4'h0;
    SS9[41][7] = 4'h0;
    SS9[42][7] = 4'h0;
    SS9[43][7] = 4'h0;
    SS9[44][7] = 4'h0;
    SS9[45][7] = 4'h0;
    SS9[46][7] = 4'h0;
    SS9[47][7] = 4'h0;
    SS9[0][8] = 4'h0;
    SS9[1][8] = 4'h0;
    SS9[2][8] = 4'h0;
    SS9[3][8] = 4'h0;
    SS9[4][8] = 4'h0;
    SS9[5][8] = 4'h0;
    SS9[6][8] = 4'h0;
    SS9[7][8] = 4'h0;
    SS9[8][8] = 4'h0;
    SS9[9][8] = 4'h0;
    SS9[10][8] = 4'h0;
    SS9[11][8] = 4'h0;
    SS9[12][8] = 4'h0;
    SS9[13][8] = 4'h0;
    SS9[14][8] = 4'h0;
    SS9[15][8] = 4'h0;
    SS9[16][8] = 4'h0;
    SS9[17][8] = 4'h0;
    SS9[18][8] = 4'h3;
    SS9[19][8] = 4'h3;
    SS9[20][8] = 4'h3;
    SS9[21][8] = 4'hD;
    SS9[22][8] = 4'hD;
    SS9[23][8] = 4'hE;
    SS9[24][8] = 4'hE;
    SS9[25][8] = 4'hE;
    SS9[26][8] = 4'hE;
    SS9[27][8] = 4'h0;
    SS9[28][8] = 4'h0;
    SS9[29][8] = 4'h0;
    SS9[30][8] = 4'hC;
    SS9[31][8] = 4'hC;
    SS9[32][8] = 4'hC;
    SS9[33][8] = 4'hC;
    SS9[34][8] = 4'hC;
    SS9[35][8] = 4'hC;
    SS9[36][8] = 4'hC;
    SS9[37][8] = 4'hD;
    SS9[38][8] = 4'h0;
    SS9[39][8] = 4'h0;
    SS9[40][8] = 4'h0;
    SS9[41][8] = 4'h0;
    SS9[42][8] = 4'h0;
    SS9[43][8] = 4'h0;
    SS9[44][8] = 4'h0;
    SS9[45][8] = 4'h0;
    SS9[46][8] = 4'h0;
    SS9[47][8] = 4'h0;
    SS9[0][9] = 4'h0;
    SS9[1][9] = 4'h0;
    SS9[2][9] = 4'h0;
    SS9[3][9] = 4'h0;
    SS9[4][9] = 4'h0;
    SS9[5][9] = 4'h0;
    SS9[6][9] = 4'h0;
    SS9[7][9] = 4'h0;
    SS9[8][9] = 4'h0;
    SS9[9][9] = 4'h0;
    SS9[10][9] = 4'h0;
    SS9[11][9] = 4'h0;
    SS9[12][9] = 4'h0;
    SS9[13][9] = 4'h0;
    SS9[14][9] = 4'h0;
    SS9[15][9] = 4'h0;
    SS9[16][9] = 4'h0;
    SS9[17][9] = 4'h0;
    SS9[18][9] = 4'h3;
    SS9[19][9] = 4'h3;
    SS9[20][9] = 4'hD;
    SS9[21][9] = 4'hE;
    SS9[22][9] = 4'hE;
    SS9[23][9] = 4'hE;
    SS9[24][9] = 4'hE;
    SS9[25][9] = 4'hE;
    SS9[26][9] = 4'hE;
    SS9[27][9] = 4'hE;
    SS9[28][9] = 4'hC;
    SS9[29][9] = 4'hC;
    SS9[30][9] = 4'hC;
    SS9[31][9] = 4'hC;
    SS9[32][9] = 4'hC;
    SS9[33][9] = 4'hC;
    SS9[34][9] = 4'hC;
    SS9[35][9] = 4'hC;
    SS9[36][9] = 4'hE;
    SS9[37][9] = 4'h0;
    SS9[38][9] = 4'h0;
    SS9[39][9] = 4'h0;
    SS9[40][9] = 4'h0;
    SS9[41][9] = 4'h0;
    SS9[42][9] = 4'h0;
    SS9[43][9] = 4'h0;
    SS9[44][9] = 4'h0;
    SS9[45][9] = 4'h0;
    SS9[46][9] = 4'h0;
    SS9[47][9] = 4'h0;
    SS9[0][10] = 4'h0;
    SS9[1][10] = 4'h0;
    SS9[2][10] = 4'h0;
    SS9[3][10] = 4'h0;
    SS9[4][10] = 4'h0;
    SS9[5][10] = 4'h0;
    SS9[6][10] = 4'h0;
    SS9[7][10] = 4'h0;
    SS9[8][10] = 4'h0;
    SS9[9][10] = 4'h0;
    SS9[10][10] = 4'h0;
    SS9[11][10] = 4'h0;
    SS9[12][10] = 4'h0;
    SS9[13][10] = 4'h0;
    SS9[14][10] = 4'h0;
    SS9[15][10] = 4'h0;
    SS9[16][10] = 4'h0;
    SS9[17][10] = 4'h0;
    SS9[18][10] = 4'hD;
    SS9[19][10] = 4'hD;
    SS9[20][10] = 4'hD;
    SS9[21][10] = 4'hD;
    SS9[22][10] = 4'hE;
    SS9[23][10] = 4'hE;
    SS9[24][10] = 4'hE;
    SS9[25][10] = 4'hE;
    SS9[26][10] = 4'hC;
    SS9[27][10] = 4'hC;
    SS9[28][10] = 4'hC;
    SS9[29][10] = 4'hC;
    SS9[30][10] = 4'hC;
    SS9[31][10] = 4'hC;
    SS9[32][10] = 4'hC;
    SS9[33][10] = 4'hD;
    SS9[34][10] = 4'hE;
    SS9[35][10] = 4'hE;
    SS9[36][10] = 4'hE;
    SS9[37][10] = 4'hE;
    SS9[38][10] = 4'h0;
    SS9[39][10] = 4'h0;
    SS9[40][10] = 4'h0;
    SS9[41][10] = 4'h0;
    SS9[42][10] = 4'h0;
    SS9[43][10] = 4'h0;
    SS9[44][10] = 4'h0;
    SS9[45][10] = 4'h0;
    SS9[46][10] = 4'h0;
    SS9[47][10] = 4'h0;
    SS9[0][11] = 4'h0;
    SS9[1][11] = 4'h0;
    SS9[2][11] = 4'h0;
    SS9[3][11] = 4'h0;
    SS9[4][11] = 4'h0;
    SS9[5][11] = 4'h0;
    SS9[6][11] = 4'h0;
    SS9[7][11] = 4'h0;
    SS9[8][11] = 4'h0;
    SS9[9][11] = 4'h0;
    SS9[10][11] = 4'h0;
    SS9[11][11] = 4'h0;
    SS9[12][11] = 4'h0;
    SS9[13][11] = 4'h0;
    SS9[14][11] = 4'h0;
    SS9[15][11] = 4'h0;
    SS9[16][11] = 4'h0;
    SS9[17][11] = 4'h0;
    SS9[18][11] = 4'h0;
    SS9[19][11] = 4'hD;
    SS9[20][11] = 4'hD;
    SS9[21][11] = 4'hD;
    SS9[22][11] = 4'hE;
    SS9[23][11] = 4'hE;
    SS9[24][11] = 4'hE;
    SS9[25][11] = 4'hC;
    SS9[26][11] = 4'hC;
    SS9[27][11] = 4'hC;
    SS9[28][11] = 4'hC;
    SS9[29][11] = 4'hC;
    SS9[30][11] = 4'hC;
    SS9[31][11] = 4'hC;
    SS9[32][11] = 4'hD;
    SS9[33][11] = 4'hD;
    SS9[34][11] = 4'hD;
    SS9[35][11] = 4'hE;
    SS9[36][11] = 4'hE;
    SS9[37][11] = 4'hE;
    SS9[38][11] = 4'h0;
    SS9[39][11] = 4'h0;
    SS9[40][11] = 4'h0;
    SS9[41][11] = 4'h0;
    SS9[42][11] = 4'h0;
    SS9[43][11] = 4'h0;
    SS9[44][11] = 4'h0;
    SS9[45][11] = 4'h0;
    SS9[46][11] = 4'h0;
    SS9[47][11] = 4'h0;
    SS9[0][12] = 4'h0;
    SS9[1][12] = 4'h0;
    SS9[2][12] = 4'h0;
    SS9[3][12] = 4'h0;
    SS9[4][12] = 4'h0;
    SS9[5][12] = 4'h0;
    SS9[6][12] = 4'h0;
    SS9[7][12] = 4'h0;
    SS9[8][12] = 4'h0;
    SS9[9][12] = 4'h0;
    SS9[10][12] = 4'h0;
    SS9[11][12] = 4'h0;
    SS9[12][12] = 4'h0;
    SS9[13][12] = 4'h0;
    SS9[14][12] = 4'h0;
    SS9[15][12] = 4'h0;
    SS9[16][12] = 4'h0;
    SS9[17][12] = 4'h0;
    SS9[18][12] = 4'h0;
    SS9[19][12] = 4'hD;
    SS9[20][12] = 4'hD;
    SS9[21][12] = 4'hD;
    SS9[22][12] = 4'hE;
    SS9[23][12] = 4'hE;
    SS9[24][12] = 4'hE;
    SS9[25][12] = 4'hE;
    SS9[26][12] = 4'hC;
    SS9[27][12] = 4'hC;
    SS9[28][12] = 4'hC;
    SS9[29][12] = 4'hC;
    SS9[30][12] = 4'hC;
    SS9[31][12] = 4'hC;
    SS9[32][12] = 4'hD;
    SS9[33][12] = 4'hD;
    SS9[34][12] = 4'hD;
    SS9[35][12] = 4'hE;
    SS9[36][12] = 4'h0;
    SS9[37][12] = 4'h0;
    SS9[38][12] = 4'h0;
    SS9[39][12] = 4'h0;
    SS9[40][12] = 4'h0;
    SS9[41][12] = 4'h0;
    SS9[42][12] = 4'h0;
    SS9[43][12] = 4'h0;
    SS9[44][12] = 4'h0;
    SS9[45][12] = 4'h0;
    SS9[46][12] = 4'h0;
    SS9[47][12] = 4'h0;
    SS9[0][13] = 4'h0;
    SS9[1][13] = 4'h0;
    SS9[2][13] = 4'h0;
    SS9[3][13] = 4'h0;
    SS9[4][13] = 4'h0;
    SS9[5][13] = 4'h0;
    SS9[6][13] = 4'h0;
    SS9[7][13] = 4'h0;
    SS9[8][13] = 4'h0;
    SS9[9][13] = 4'h0;
    SS9[10][13] = 4'h0;
    SS9[11][13] = 4'h0;
    SS9[12][13] = 4'h0;
    SS9[13][13] = 4'h0;
    SS9[14][13] = 4'h0;
    SS9[15][13] = 4'h0;
    SS9[16][13] = 4'h0;
    SS9[17][13] = 4'h0;
    SS9[18][13] = 4'hD;
    SS9[19][13] = 4'hD;
    SS9[20][13] = 4'hD;
    SS9[21][13] = 4'hD;
    SS9[22][13] = 4'hD;
    SS9[23][13] = 4'hE;
    SS9[24][13] = 4'hE;
    SS9[25][13] = 4'hE;
    SS9[26][13] = 4'hC;
    SS9[27][13] = 4'hC;
    SS9[28][13] = 4'hC;
    SS9[29][13] = 4'hC;
    SS9[30][13] = 4'hC;
    SS9[31][13] = 4'hC;
    SS9[32][13] = 4'hD;
    SS9[33][13] = 4'hD;
    SS9[34][13] = 4'hE;
    SS9[35][13] = 4'hE;
    SS9[36][13] = 4'h0;
    SS9[37][13] = 4'h0;
    SS9[38][13] = 4'h0;
    SS9[39][13] = 4'h0;
    SS9[40][13] = 4'h0;
    SS9[41][13] = 4'h0;
    SS9[42][13] = 4'h0;
    SS9[43][13] = 4'h0;
    SS9[44][13] = 4'h0;
    SS9[45][13] = 4'h0;
    SS9[46][13] = 4'h0;
    SS9[47][13] = 4'h0;
    SS9[0][14] = 4'h0;
    SS9[1][14] = 4'h0;
    SS9[2][14] = 4'h0;
    SS9[3][14] = 4'h0;
    SS9[4][14] = 4'h0;
    SS9[5][14] = 4'h0;
    SS9[6][14] = 4'h0;
    SS9[7][14] = 4'h0;
    SS9[8][14] = 4'h0;
    SS9[9][14] = 4'h0;
    SS9[10][14] = 4'h0;
    SS9[11][14] = 4'h0;
    SS9[12][14] = 4'h0;
    SS9[13][14] = 4'h0;
    SS9[14][14] = 4'h0;
    SS9[15][14] = 4'h0;
    SS9[16][14] = 4'h3;
    SS9[17][14] = 4'hD;
    SS9[18][14] = 4'hD;
    SS9[19][14] = 4'hD;
    SS9[20][14] = 4'hD;
    SS9[21][14] = 4'hD;
    SS9[22][14] = 4'hD;
    SS9[23][14] = 4'hE;
    SS9[24][14] = 4'hC;
    SS9[25][14] = 4'hC;
    SS9[26][14] = 4'hC;
    SS9[27][14] = 4'hC;
    SS9[28][14] = 4'hC;
    SS9[29][14] = 4'hC;
    SS9[30][14] = 4'hC;
    SS9[31][14] = 4'hD;
    SS9[32][14] = 4'hD;
    SS9[33][14] = 4'hE;
    SS9[34][14] = 4'hE;
    SS9[35][14] = 4'hE;
    SS9[36][14] = 4'h0;
    SS9[37][14] = 4'h0;
    SS9[38][14] = 4'h0;
    SS9[39][14] = 4'h0;
    SS9[40][14] = 4'h0;
    SS9[41][14] = 4'h0;
    SS9[42][14] = 4'h0;
    SS9[43][14] = 4'h0;
    SS9[44][14] = 4'h0;
    SS9[45][14] = 4'h0;
    SS9[46][14] = 4'h0;
    SS9[47][14] = 4'h0;
    SS9[0][15] = 4'h0;
    SS9[1][15] = 4'h0;
    SS9[2][15] = 4'h0;
    SS9[3][15] = 4'h0;
    SS9[4][15] = 4'h0;
    SS9[5][15] = 4'h0;
    SS9[6][15] = 4'h0;
    SS9[7][15] = 4'h0;
    SS9[8][15] = 4'h0;
    SS9[9][15] = 4'h0;
    SS9[10][15] = 4'h0;
    SS9[11][15] = 4'h0;
    SS9[12][15] = 4'h0;
    SS9[13][15] = 4'h0;
    SS9[14][15] = 4'h3;
    SS9[15][15] = 4'h3;
    SS9[16][15] = 4'h3;
    SS9[17][15] = 4'hD;
    SS9[18][15] = 4'hD;
    SS9[19][15] = 4'hD;
    SS9[20][15] = 4'hD;
    SS9[21][15] = 4'hE;
    SS9[22][15] = 4'hE;
    SS9[23][15] = 4'hE;
    SS9[24][15] = 4'hC;
    SS9[25][15] = 4'hC;
    SS9[26][15] = 4'hC;
    SS9[27][15] = 4'hC;
    SS9[28][15] = 4'hC;
    SS9[29][15] = 4'hC;
    SS9[30][15] = 4'hD;
    SS9[31][15] = 4'hD;
    SS9[32][15] = 4'hD;
    SS9[33][15] = 4'hE;
    SS9[34][15] = 4'hE;
    SS9[35][15] = 4'hE;
    SS9[36][15] = 4'hE;
    SS9[37][15] = 4'h0;
    SS9[38][15] = 4'h0;
    SS9[39][15] = 4'h0;
    SS9[40][15] = 4'h0;
    SS9[41][15] = 4'h0;
    SS9[42][15] = 4'h0;
    SS9[43][15] = 4'h0;
    SS9[44][15] = 4'h0;
    SS9[45][15] = 4'h0;
    SS9[46][15] = 4'h0;
    SS9[47][15] = 4'h0;
    SS9[0][16] = 4'h0;
    SS9[1][16] = 4'h0;
    SS9[2][16] = 4'h0;
    SS9[3][16] = 4'h0;
    SS9[4][16] = 4'h0;
    SS9[5][16] = 4'h0;
    SS9[6][16] = 4'h0;
    SS9[7][16] = 4'h0;
    SS9[8][16] = 4'h0;
    SS9[9][16] = 4'h0;
    SS9[10][16] = 4'h0;
    SS9[11][16] = 4'h0;
    SS9[12][16] = 4'h0;
    SS9[13][16] = 4'h0;
    SS9[14][16] = 4'h3;
    SS9[15][16] = 4'h3;
    SS9[16][16] = 4'h3;
    SS9[17][16] = 4'h3;
    SS9[18][16] = 4'hD;
    SS9[19][16] = 4'hD;
    SS9[20][16] = 4'hD;
    SS9[21][16] = 4'hE;
    SS9[22][16] = 4'hE;
    SS9[23][16] = 4'hE;
    SS9[24][16] = 4'hC;
    SS9[25][16] = 4'hC;
    SS9[26][16] = 4'hC;
    SS9[27][16] = 4'hC;
    SS9[28][16] = 4'hC;
    SS9[29][16] = 4'hC;
    SS9[30][16] = 4'hC;
    SS9[31][16] = 4'hD;
    SS9[32][16] = 4'hD;
    SS9[33][16] = 4'hD;
    SS9[34][16] = 4'h0;
    SS9[35][16] = 4'h0;
    SS9[36][16] = 4'h0;
    SS9[37][16] = 4'h0;
    SS9[38][16] = 4'h0;
    SS9[39][16] = 4'h0;
    SS9[40][16] = 4'h0;
    SS9[41][16] = 4'h0;
    SS9[42][16] = 4'h0;
    SS9[43][16] = 4'h0;
    SS9[44][16] = 4'h0;
    SS9[45][16] = 4'h0;
    SS9[46][16] = 4'h0;
    SS9[47][16] = 4'h0;
    SS9[0][17] = 4'h0;
    SS9[1][17] = 4'h0;
    SS9[2][17] = 4'h0;
    SS9[3][17] = 4'h0;
    SS9[4][17] = 4'h0;
    SS9[5][17] = 4'h0;
    SS9[6][17] = 4'h0;
    SS9[7][17] = 4'h0;
    SS9[8][17] = 4'h0;
    SS9[9][17] = 4'h0;
    SS9[10][17] = 4'h0;
    SS9[11][17] = 4'h0;
    SS9[12][17] = 4'h0;
    SS9[13][17] = 4'h0;
    SS9[14][17] = 4'h0;
    SS9[15][17] = 4'h3;
    SS9[16][17] = 4'hD;
    SS9[17][17] = 4'hD;
    SS9[18][17] = 4'hD;
    SS9[19][17] = 4'hD;
    SS9[20][17] = 4'hD;
    SS9[21][17] = 4'hE;
    SS9[22][17] = 4'hE;
    SS9[23][17] = 4'hE;
    SS9[24][17] = 4'hC;
    SS9[25][17] = 4'hC;
    SS9[26][17] = 4'hC;
    SS9[27][17] = 4'hC;
    SS9[28][17] = 4'hC;
    SS9[29][17] = 4'hC;
    SS9[30][17] = 4'hC;
    SS9[31][17] = 4'hD;
    SS9[32][17] = 4'hE;
    SS9[33][17] = 4'hE;
    SS9[34][17] = 4'h0;
    SS9[35][17] = 4'h0;
    SS9[36][17] = 4'h0;
    SS9[37][17] = 4'h0;
    SS9[38][17] = 4'h0;
    SS9[39][17] = 4'h0;
    SS9[40][17] = 4'h0;
    SS9[41][17] = 4'h0;
    SS9[42][17] = 4'h0;
    SS9[43][17] = 4'h0;
    SS9[44][17] = 4'h0;
    SS9[45][17] = 4'h0;
    SS9[46][17] = 4'h0;
    SS9[47][17] = 4'h0;
    SS9[0][18] = 4'h0;
    SS9[1][18] = 4'h0;
    SS9[2][18] = 4'h0;
    SS9[3][18] = 4'h0;
    SS9[4][18] = 4'h0;
    SS9[5][18] = 4'h0;
    SS9[6][18] = 4'h0;
    SS9[7][18] = 4'h0;
    SS9[8][18] = 4'h0;
    SS9[9][18] = 4'h0;
    SS9[10][18] = 4'h0;
    SS9[11][18] = 4'h0;
    SS9[12][18] = 4'h0;
    SS9[13][18] = 4'h0;
    SS9[14][18] = 4'h0;
    SS9[15][18] = 4'hD;
    SS9[16][18] = 4'hD;
    SS9[17][18] = 4'hD;
    SS9[18][18] = 4'hD;
    SS9[19][18] = 4'hD;
    SS9[20][18] = 4'hD;
    SS9[21][18] = 4'hD;
    SS9[22][18] = 4'hC;
    SS9[23][18] = 4'hC;
    SS9[24][18] = 4'hC;
    SS9[25][18] = 4'hC;
    SS9[26][18] = 4'hC;
    SS9[27][18] = 4'hC;
    SS9[28][18] = 4'hC;
    SS9[29][18] = 4'hC;
    SS9[30][18] = 4'hE;
    SS9[31][18] = 4'hE;
    SS9[32][18] = 4'hE;
    SS9[33][18] = 4'hE;
    SS9[34][18] = 4'hE;
    SS9[35][18] = 4'h0;
    SS9[36][18] = 4'h0;
    SS9[37][18] = 4'h0;
    SS9[38][18] = 4'h0;
    SS9[39][18] = 4'h0;
    SS9[40][18] = 4'h0;
    SS9[41][18] = 4'h0;
    SS9[42][18] = 4'h0;
    SS9[43][18] = 4'h0;
    SS9[44][18] = 4'h0;
    SS9[45][18] = 4'h0;
    SS9[46][18] = 4'h0;
    SS9[47][18] = 4'h0;
    SS9[0][19] = 4'h0;
    SS9[1][19] = 4'h0;
    SS9[2][19] = 4'h0;
    SS9[3][19] = 4'h0;
    SS9[4][19] = 4'h0;
    SS9[5][19] = 4'h0;
    SS9[6][19] = 4'h0;
    SS9[7][19] = 4'h0;
    SS9[8][19] = 4'h0;
    SS9[9][19] = 4'h0;
    SS9[10][19] = 4'h0;
    SS9[11][19] = 4'h0;
    SS9[12][19] = 4'h0;
    SS9[13][19] = 4'h0;
    SS9[14][19] = 4'h0;
    SS9[15][19] = 4'h0;
    SS9[16][19] = 4'hD;
    SS9[17][19] = 4'hD;
    SS9[18][19] = 4'hD;
    SS9[19][19] = 4'hC;
    SS9[20][19] = 4'hC;
    SS9[21][19] = 4'hC;
    SS9[22][19] = 4'hC;
    SS9[23][19] = 4'hC;
    SS9[24][19] = 4'hC;
    SS9[25][19] = 4'hC;
    SS9[26][19] = 4'hC;
    SS9[27][19] = 4'hD;
    SS9[28][19] = 4'hD;
    SS9[29][19] = 4'hE;
    SS9[30][19] = 4'hE;
    SS9[31][19] = 4'hE;
    SS9[32][19] = 4'hE;
    SS9[33][19] = 4'hE;
    SS9[34][19] = 4'hE;
    SS9[35][19] = 4'h0;
    SS9[36][19] = 4'h0;
    SS9[37][19] = 4'h0;
    SS9[38][19] = 4'h0;
    SS9[39][19] = 4'h0;
    SS9[40][19] = 4'h0;
    SS9[41][19] = 4'h0;
    SS9[42][19] = 4'h0;
    SS9[43][19] = 4'h0;
    SS9[44][19] = 4'h0;
    SS9[45][19] = 4'h0;
    SS9[46][19] = 4'h0;
    SS9[47][19] = 4'h0;
    SS9[0][20] = 4'h0;
    SS9[1][20] = 4'h0;
    SS9[2][20] = 4'h0;
    SS9[3][20] = 4'h0;
    SS9[4][20] = 4'h0;
    SS9[5][20] = 4'h0;
    SS9[6][20] = 4'h0;
    SS9[7][20] = 4'h0;
    SS9[8][20] = 4'h0;
    SS9[9][20] = 4'h0;
    SS9[10][20] = 4'h0;
    SS9[11][20] = 4'h0;
    SS9[12][20] = 4'h0;
    SS9[13][20] = 4'h0;
    SS9[14][20] = 4'h0;
    SS9[15][20] = 4'h0;
    SS9[16][20] = 4'hD;
    SS9[17][20] = 4'hD;
    SS9[18][20] = 4'hD;
    SS9[19][20] = 4'hC;
    SS9[20][20] = 4'hC;
    SS9[21][20] = 4'hC;
    SS9[22][20] = 4'hC;
    SS9[23][20] = 4'hC;
    SS9[24][20] = 4'hC;
    SS9[25][20] = 4'hC;
    SS9[26][20] = 4'hD;
    SS9[27][20] = 4'hD;
    SS9[28][20] = 4'hD;
    SS9[29][20] = 4'hE;
    SS9[30][20] = 4'hE;
    SS9[31][20] = 4'hE;
    SS9[32][20] = 4'hE;
    SS9[33][20] = 4'hE;
    SS9[34][20] = 4'hE;
    SS9[35][20] = 4'h0;
    SS9[36][20] = 4'h0;
    SS9[37][20] = 4'h0;
    SS9[38][20] = 4'h0;
    SS9[39][20] = 4'h0;
    SS9[40][20] = 4'h0;
    SS9[41][20] = 4'h0;
    SS9[42][20] = 4'h0;
    SS9[43][20] = 4'h0;
    SS9[44][20] = 4'h0;
    SS9[45][20] = 4'h0;
    SS9[46][20] = 4'h0;
    SS9[47][20] = 4'h0;
    SS9[0][21] = 4'h0;
    SS9[1][21] = 4'h0;
    SS9[2][21] = 4'h0;
    SS9[3][21] = 4'h0;
    SS9[4][21] = 4'h0;
    SS9[5][21] = 4'h0;
    SS9[6][21] = 4'h0;
    SS9[7][21] = 4'h0;
    SS9[8][21] = 4'h0;
    SS9[9][21] = 4'h0;
    SS9[10][21] = 4'h0;
    SS9[11][21] = 4'h0;
    SS9[12][21] = 4'h0;
    SS9[13][21] = 4'h0;
    SS9[14][21] = 4'hE;
    SS9[15][21] = 4'hC;
    SS9[16][21] = 4'hC;
    SS9[17][21] = 4'hD;
    SS9[18][21] = 4'hD;
    SS9[19][21] = 4'hD;
    SS9[20][21] = 4'hC;
    SS9[21][21] = 4'hC;
    SS9[22][21] = 4'hD;
    SS9[23][21] = 4'hC;
    SS9[24][21] = 4'hC;
    SS9[25][21] = 4'hC;
    SS9[26][21] = 4'hD;
    SS9[27][21] = 4'hD;
    SS9[28][21] = 4'hD;
    SS9[29][21] = 4'hE;
    SS9[30][21] = 4'hE;
    SS9[31][21] = 4'hE;
    SS9[32][21] = 4'hE;
    SS9[33][21] = 4'hE;
    SS9[34][21] = 4'hE;
    SS9[35][21] = 4'hE;
    SS9[36][21] = 4'h0;
    SS9[37][21] = 4'h0;
    SS9[38][21] = 4'hE;
    SS9[39][21] = 4'h0;
    SS9[40][21] = 4'h0;
    SS9[41][21] = 4'h0;
    SS9[42][21] = 4'h0;
    SS9[43][21] = 4'h0;
    SS9[44][21] = 4'h0;
    SS9[45][21] = 4'h0;
    SS9[46][21] = 4'h0;
    SS9[47][21] = 4'h0;
    SS9[0][22] = 4'h0;
    SS9[1][22] = 4'h0;
    SS9[2][22] = 4'h0;
    SS9[3][22] = 4'h0;
    SS9[4][22] = 4'h0;
    SS9[5][22] = 4'h0;
    SS9[6][22] = 4'h0;
    SS9[7][22] = 4'h0;
    SS9[8][22] = 4'h0;
    SS9[9][22] = 4'h0;
    SS9[10][22] = 4'h0;
    SS9[11][22] = 4'h0;
    SS9[12][22] = 4'hD;
    SS9[13][22] = 4'hD;
    SS9[14][22] = 4'hC;
    SS9[15][22] = 4'hC;
    SS9[16][22] = 4'hC;
    SS9[17][22] = 4'hD;
    SS9[18][22] = 4'hD;
    SS9[19][22] = 4'hD;
    SS9[20][22] = 4'hD;
    SS9[21][22] = 4'hD;
    SS9[22][22] = 4'hD;
    SS9[23][22] = 4'hC;
    SS9[24][22] = 4'hC;
    SS9[25][22] = 4'hC;
    SS9[26][22] = 4'hC;
    SS9[27][22] = 4'hD;
    SS9[28][22] = 4'hD;
    SS9[29][22] = 4'hD;
    SS9[30][22] = 4'hE;
    SS9[31][22] = 4'hE;
    SS9[32][22] = 4'hE;
    SS9[33][22] = 4'hE;
    SS9[34][22] = 4'hE;
    SS9[35][22] = 4'hD;
    SS9[36][22] = 4'hE;
    SS9[37][22] = 4'hE;
    SS9[38][22] = 4'hE;
    SS9[39][22] = 4'h0;
    SS9[40][22] = 4'h0;
    SS9[41][22] = 4'h0;
    SS9[42][22] = 4'h0;
    SS9[43][22] = 4'h0;
    SS9[44][22] = 4'h0;
    SS9[45][22] = 4'h0;
    SS9[46][22] = 4'h0;
    SS9[47][22] = 4'h0;
    SS9[0][23] = 4'h0;
    SS9[1][23] = 4'h0;
    SS9[2][23] = 4'h0;
    SS9[3][23] = 4'h0;
    SS9[4][23] = 4'h0;
    SS9[5][23] = 4'h0;
    SS9[6][23] = 4'h0;
    SS9[7][23] = 4'h0;
    SS9[8][23] = 4'h0;
    SS9[9][23] = 4'h0;
    SS9[10][23] = 4'hD;
    SS9[11][23] = 4'hD;
    SS9[12][23] = 4'hD;
    SS9[13][23] = 4'hD;
    SS9[14][23] = 4'hC;
    SS9[15][23] = 4'hC;
    SS9[16][23] = 4'hC;
    SS9[17][23] = 4'hA;
    SS9[18][23] = 4'hA;
    SS9[19][23] = 4'hA;
    SS9[20][23] = 4'hA;
    SS9[21][23] = 4'hD;
    SS9[22][23] = 4'hD;
    SS9[23][23] = 4'hD;
    SS9[24][23] = 4'hC;
    SS9[25][23] = 4'hC;
    SS9[26][23] = 4'hC;
    SS9[27][23] = 4'hD;
    SS9[28][23] = 4'hD;
    SS9[29][23] = 4'hD;
    SS9[30][23] = 4'hE;
    SS9[31][23] = 4'hE;
    SS9[32][23] = 4'hE;
    SS9[33][23] = 4'hD;
    SS9[34][23] = 4'hD;
    SS9[35][23] = 4'hD;
    SS9[36][23] = 4'hD;
    SS9[37][23] = 4'hE;
    SS9[38][23] = 4'hE;
    SS9[39][23] = 4'hE;
    SS9[40][23] = 4'h0;
    SS9[41][23] = 4'hE;
    SS9[42][23] = 4'hE;
    SS9[43][23] = 4'h0;
    SS9[44][23] = 4'h0;
    SS9[45][23] = 4'h0;
    SS9[46][23] = 4'h0;
    SS9[47][23] = 4'h0;
    SS9[0][24] = 4'h0;
    SS9[1][24] = 4'h0;
    SS9[2][24] = 4'h0;
    SS9[3][24] = 4'h0;
    SS9[4][24] = 4'h0;
    SS9[5][24] = 4'h0;
    SS9[6][24] = 4'h0;
    SS9[7][24] = 4'hD;
    SS9[8][24] = 4'hD;
    SS9[9][24] = 4'hD;
    SS9[10][24] = 4'hD;
    SS9[11][24] = 4'hD;
    SS9[12][24] = 4'hD;
    SS9[13][24] = 4'hD;
    SS9[14][24] = 4'hD;
    SS9[15][24] = 4'hC;
    SS9[16][24] = 4'hC;
    SS9[17][24] = 4'hC;
    SS9[18][24] = 4'hA;
    SS9[19][24] = 4'hA;
    SS9[20][24] = 4'hA;
    SS9[21][24] = 4'hD;
    SS9[22][24] = 4'hD;
    SS9[23][24] = 4'hD;
    SS9[24][24] = 4'hC;
    SS9[25][24] = 4'hC;
    SS9[26][24] = 4'hC;
    SS9[27][24] = 4'hD;
    SS9[28][24] = 4'hD;
    SS9[29][24] = 4'hD;
    SS9[30][24] = 4'hD;
    SS9[31][24] = 4'hC;
    SS9[32][24] = 4'hC;
    SS9[33][24] = 4'hC;
    SS9[34][24] = 4'hD;
    SS9[35][24] = 4'hD;
    SS9[36][24] = 4'hD;
    SS9[37][24] = 4'hE;
    SS9[38][24] = 4'hD;
    SS9[39][24] = 4'hD;
    SS9[40][24] = 4'hE;
    SS9[41][24] = 4'hE;
    SS9[42][24] = 4'hE;
    SS9[43][24] = 4'h0;
    SS9[44][24] = 4'h0;
    SS9[45][24] = 4'h0;
    SS9[46][24] = 4'hD;
    SS9[47][24] = 4'h0;
    SS9[0][25] = 4'h0;
    SS9[1][25] = 4'h0;
    SS9[2][25] = 4'h0;
    SS9[3][25] = 4'h0;
    SS9[4][25] = 4'h0;
    SS9[5][25] = 4'hD;
    SS9[6][25] = 4'hD;
    SS9[7][25] = 4'hD;
    SS9[8][25] = 4'hD;
    SS9[9][25] = 4'hD;
    SS9[10][25] = 4'hD;
    SS9[11][25] = 4'hD;
    SS9[12][25] = 4'hD;
    SS9[13][25] = 4'hC;
    SS9[14][25] = 4'hC;
    SS9[15][25] = 4'hC;
    SS9[16][25] = 4'hC;
    SS9[17][25] = 4'hC;
    SS9[18][25] = 4'hA;
    SS9[19][25] = 4'hA;
    SS9[20][25] = 4'hA;
    SS9[21][25] = 4'hD;
    SS9[22][25] = 4'hD;
    SS9[23][25] = 4'hD;
    SS9[24][25] = 4'hD;
    SS9[25][25] = 4'hC;
    SS9[26][25] = 4'hC;
    SS9[27][25] = 4'hC;
    SS9[28][25] = 4'hC;
    SS9[29][25] = 4'hC;
    SS9[30][25] = 4'hC;
    SS9[31][25] = 4'hC;
    SS9[32][25] = 4'hC;
    SS9[33][25] = 4'hC;
    SS9[34][25] = 4'hD;
    SS9[35][25] = 4'hD;
    SS9[36][25] = 4'hC;
    SS9[37][25] = 4'hD;
    SS9[38][25] = 4'hD;
    SS9[39][25] = 4'hD;
    SS9[40][25] = 4'hD;
    SS9[41][25] = 4'hE;
    SS9[42][25] = 4'hE;
    SS9[43][25] = 4'hE;
    SS9[44][25] = 4'hD;
    SS9[45][25] = 4'hD;
    SS9[46][25] = 4'hD;
    SS9[47][25] = 4'h0;
    SS9[0][26] = 4'h0;
    SS9[1][26] = 4'h0;
    SS9[2][26] = 4'h0;
    SS9[3][26] = 4'h0;
    SS9[4][26] = 4'h0;
    SS9[5][26] = 4'h0;
    SS9[6][26] = 4'hD;
    SS9[7][26] = 4'hD;
    SS9[8][26] = 4'hD;
    SS9[9][26] = 4'hD;
    SS9[10][26] = 4'hC;
    SS9[11][26] = 4'hC;
    SS9[12][26] = 4'hC;
    SS9[13][26] = 4'hC;
    SS9[14][26] = 4'hC;
    SS9[15][26] = 4'hC;
    SS9[16][26] = 4'hC;
    SS9[17][26] = 4'hC;
    SS9[18][26] = 4'hC;
    SS9[19][26] = 4'hA;
    SS9[20][26] = 4'hA;
    SS9[21][26] = 4'hA;
    SS9[22][26] = 4'hD;
    SS9[23][26] = 4'hD;
    SS9[24][26] = 4'hD;
    SS9[25][26] = 4'hC;
    SS9[26][26] = 4'hC;
    SS9[27][26] = 4'hC;
    SS9[28][26] = 4'hC;
    SS9[29][26] = 4'hC;
    SS9[30][26] = 4'hC;
    SS9[31][26] = 4'hC;
    SS9[32][26] = 4'hC;
    SS9[33][26] = 4'hC;
    SS9[34][26] = 4'hC;
    SS9[35][26] = 4'hC;
    SS9[36][26] = 4'hC;
    SS9[37][26] = 4'hC;
    SS9[38][26] = 4'hD;
    SS9[39][26] = 4'hD;
    SS9[40][26] = 4'hD;
    SS9[41][26] = 4'hC;
    SS9[42][26] = 4'hC;
    SS9[43][26] = 4'hC;
    SS9[44][26] = 4'hD;
    SS9[45][26] = 4'hD;
    SS9[46][26] = 4'hD;
    SS9[47][26] = 4'h0;
    SS9[0][27] = 4'h0;
    SS9[1][27] = 4'h0;
    SS9[2][27] = 4'h0;
    SS9[3][27] = 4'h0;
    SS9[4][27] = 4'h0;
    SS9[5][27] = 4'h0;
    SS9[6][27] = 4'hD;
    SS9[7][27] = 4'hD;
    SS9[8][27] = 4'hC;
    SS9[9][27] = 4'hC;
    SS9[10][27] = 4'hC;
    SS9[11][27] = 4'hC;
    SS9[12][27] = 4'hC;
    SS9[13][27] = 4'hC;
    SS9[14][27] = 4'hC;
    SS9[15][27] = 4'hC;
    SS9[16][27] = 4'hC;
    SS9[17][27] = 4'hC;
    SS9[18][27] = 4'hC;
    SS9[19][27] = 4'hA;
    SS9[20][27] = 4'hA;
    SS9[21][27] = 4'hA;
    SS9[22][27] = 4'hD;
    SS9[23][27] = 4'hC;
    SS9[24][27] = 4'hC;
    SS9[25][27] = 4'hC;
    SS9[26][27] = 4'hC;
    SS9[27][27] = 4'hC;
    SS9[28][27] = 4'hC;
    SS9[29][27] = 4'hC;
    SS9[30][27] = 4'hC;
    SS9[31][27] = 4'hC;
    SS9[32][27] = 4'hC;
    SS9[33][27] = 4'hC;
    SS9[34][27] = 4'hC;
    SS9[35][27] = 4'hC;
    SS9[36][27] = 4'hC;
    SS9[37][27] = 4'hC;
    SS9[38][27] = 4'hD;
    SS9[39][27] = 4'hC;
    SS9[40][27] = 4'hC;
    SS9[41][27] = 4'hC;
    SS9[42][27] = 4'hC;
    SS9[43][27] = 4'hC;
    SS9[44][27] = 4'hC;
    SS9[45][27] = 4'hD;
    SS9[46][27] = 4'hD;
    SS9[47][27] = 4'hC;
    SS9[0][28] = 4'h0;
    SS9[1][28] = 4'h0;
    SS9[2][28] = 4'h0;
    SS9[3][28] = 4'h0;
    SS9[4][28] = 4'h0;
    SS9[5][28] = 4'hC;
    SS9[6][28] = 4'hC;
    SS9[7][28] = 4'hC;
    SS9[8][28] = 4'hC;
    SS9[9][28] = 4'hC;
    SS9[10][28] = 4'hC;
    SS9[11][28] = 4'hC;
    SS9[12][28] = 4'hC;
    SS9[13][28] = 4'hC;
    SS9[14][28] = 4'hC;
    SS9[15][28] = 4'hC;
    SS9[16][28] = 4'hC;
    SS9[17][28] = 4'hC;
    SS9[18][28] = 4'hC;
    SS9[19][28] = 4'hA;
    SS9[20][28] = 4'hA;
    SS9[21][28] = 4'hD;
    SS9[22][28] = 4'hD;
    SS9[23][28] = 4'hC;
    SS9[24][28] = 4'hC;
    SS9[25][28] = 4'hC;
    SS9[26][28] = 4'hC;
    SS9[27][28] = 4'hC;
    SS9[28][28] = 4'hC;
    SS9[29][28] = 4'hC;
    SS9[30][28] = 4'hC;
    SS9[31][28] = 4'hC;
    SS9[32][28] = 4'hC;
    SS9[33][28] = 4'hC;
    SS9[34][28] = 4'hC;
    SS9[35][28] = 4'hC;
    SS9[36][28] = 4'hC;
    SS9[37][28] = 4'hC;
    SS9[38][28] = 4'hC;
    SS9[39][28] = 4'hC;
    SS9[40][28] = 4'hC;
    SS9[41][28] = 4'hC;
    SS9[42][28] = 4'hC;
    SS9[43][28] = 4'hC;
    SS9[44][28] = 4'hC;
    SS9[45][28] = 4'hC;
    SS9[46][28] = 4'hC;
    SS9[47][28] = 4'hC;
    SS9[0][29] = 4'h0;
    SS9[1][29] = 4'h0;
    SS9[2][29] = 4'h0;
    SS9[3][29] = 4'hC;
    SS9[4][29] = 4'hC;
    SS9[5][29] = 4'hC;
    SS9[6][29] = 4'hC;
    SS9[7][29] = 4'hC;
    SS9[8][29] = 4'hC;
    SS9[9][29] = 4'hC;
    SS9[10][29] = 4'hC;
    SS9[11][29] = 4'hC;
    SS9[12][29] = 4'hC;
    SS9[13][29] = 4'hC;
    SS9[14][29] = 4'hC;
    SS9[15][29] = 4'hC;
    SS9[16][29] = 4'hC;
    SS9[17][29] = 4'hC;
    SS9[18][29] = 4'hC;
    SS9[19][29] = 4'hC;
    SS9[20][29] = 4'hD;
    SS9[21][29] = 4'hD;
    SS9[22][29] = 4'hD;
    SS9[23][29] = 4'hC;
    SS9[24][29] = 4'hC;
    SS9[25][29] = 4'hC;
    SS9[26][29] = 4'hE;
    SS9[27][29] = 4'hE;
    SS9[28][29] = 4'hE;
    SS9[29][29] = 4'hC;
    SS9[30][29] = 4'hC;
    SS9[31][29] = 4'hC;
    SS9[32][29] = 4'hC;
    SS9[33][29] = 4'hC;
    SS9[34][29] = 4'hC;
    SS9[35][29] = 4'hC;
    SS9[36][29] = 4'hC;
    SS9[37][29] = 4'hC;
    SS9[38][29] = 4'hC;
    SS9[39][29] = 4'hC;
    SS9[40][29] = 4'hC;
    SS9[41][29] = 4'hC;
    SS9[42][29] = 4'hC;
    SS9[43][29] = 4'hC;
    SS9[44][29] = 4'hC;
    SS9[45][29] = 4'hC;
    SS9[46][29] = 4'hC;
    SS9[47][29] = 4'hC;
    SS9[0][30] = 4'h0;
    SS9[1][30] = 4'hC;
    SS9[2][30] = 4'hC;
    SS9[3][30] = 4'hC;
    SS9[4][30] = 4'hC;
    SS9[5][30] = 4'hC;
    SS9[6][30] = 4'hC;
    SS9[7][30] = 4'hC;
    SS9[8][30] = 4'hC;
    SS9[9][30] = 4'hC;
    SS9[10][30] = 4'hC;
    SS9[11][30] = 4'hC;
    SS9[12][30] = 4'hC;
    SS9[13][30] = 4'hC;
    SS9[14][30] = 4'hC;
    SS9[15][30] = 4'hC;
    SS9[16][30] = 4'hD;
    SS9[17][30] = 4'hC;
    SS9[18][30] = 4'hC;
    SS9[19][30] = 4'hC;
    SS9[20][30] = 4'hD;
    SS9[21][30] = 4'hD;
    SS9[22][30] = 4'hD;
    SS9[23][30] = 4'hC;
    SS9[24][30] = 4'hD;
    SS9[25][30] = 4'hD;
    SS9[26][30] = 4'hD;
    SS9[27][30] = 4'hE;
    SS9[28][30] = 4'hE;
    SS9[29][30] = 4'hE;
    SS9[30][30] = 4'hC;
    SS9[31][30] = 4'hC;
    SS9[32][30] = 4'hE;
    SS9[33][30] = 4'hC;
    SS9[34][30] = 4'hC;
    SS9[35][30] = 4'hC;
    SS9[36][30] = 4'hC;
    SS9[37][30] = 4'hC;
    SS9[38][30] = 4'hC;
    SS9[39][30] = 4'h0;
    SS9[40][30] = 4'h0;
    SS9[41][30] = 4'h0;
    SS9[42][30] = 4'h0;
    SS9[43][30] = 4'hC;
    SS9[44][30] = 4'hC;
    SS9[45][30] = 4'hC;
    SS9[46][30] = 4'hC;
    SS9[47][30] = 4'h0;
    SS9[0][31] = 4'h0;
    SS9[1][31] = 4'hC;
    SS9[2][31] = 4'hC;
    SS9[3][31] = 4'hC;
    SS9[4][31] = 4'hC;
    SS9[5][31] = 4'hC;
    SS9[6][31] = 4'hC;
    SS9[7][31] = 4'hC;
    SS9[8][31] = 4'hC;
    SS9[9][31] = 4'hC;
    SS9[10][31] = 4'hC;
    SS9[11][31] = 4'hC;
    SS9[12][31] = 4'hC;
    SS9[13][31] = 4'hC;
    SS9[14][31] = 4'hD;
    SS9[15][31] = 4'hD;
    SS9[16][31] = 4'hD;
    SS9[17][31] = 4'hC;
    SS9[18][31] = 4'hC;
    SS9[19][31] = 4'hC;
    SS9[20][31] = 4'hC;
    SS9[21][31] = 4'hD;
    SS9[22][31] = 4'hD;
    SS9[23][31] = 4'hD;
    SS9[24][31] = 4'hD;
    SS9[25][31] = 4'hD;
    SS9[26][31] = 4'hD;
    SS9[27][31] = 4'hE;
    SS9[28][31] = 4'hE;
    SS9[29][31] = 4'hD;
    SS9[30][31] = 4'hE;
    SS9[31][31] = 4'hE;
    SS9[32][31] = 4'hE;
    SS9[33][31] = 4'hE;
    SS9[34][31] = 4'hC;
    SS9[35][31] = 4'hC;
    SS9[36][31] = 4'hC;
    SS9[37][31] = 4'h0;
    SS9[38][31] = 4'h0;
    SS9[39][31] = 4'h0;
    SS9[40][31] = 4'h0;
    SS9[41][31] = 4'h0;
    SS9[42][31] = 4'h0;
    SS9[43][31] = 4'hC;
    SS9[44][31] = 4'hC;
    SS9[45][31] = 4'h0;
    SS9[46][31] = 4'h0;
    SS9[47][31] = 4'h0;
    SS9[0][32] = 4'h0;
    SS9[1][32] = 4'h0;
    SS9[2][32] = 4'hC;
    SS9[3][32] = 4'hC;
    SS9[4][32] = 4'hC;
    SS9[5][32] = 4'hC;
    SS9[6][32] = 4'hC;
    SS9[7][32] = 4'hC;
    SS9[8][32] = 4'hC;
    SS9[9][32] = 4'hC;
    SS9[10][32] = 4'hC;
    SS9[11][32] = 4'hD;
    SS9[12][32] = 4'hD;
    SS9[13][32] = 4'hD;
    SS9[14][32] = 4'hD;
    SS9[15][32] = 4'hD;
    SS9[16][32] = 4'hD;
    SS9[17][32] = 4'hD;
    SS9[18][32] = 4'hC;
    SS9[19][32] = 4'h0;
    SS9[20][32] = 4'h0;
    SS9[21][32] = 4'hD;
    SS9[22][32] = 4'hD;
    SS9[23][32] = 4'hD;
    SS9[24][32] = 4'hD;
    SS9[25][32] = 4'hD;
    SS9[26][32] = 4'hD;
    SS9[27][32] = 4'hD;
    SS9[28][32] = 4'hD;
    SS9[29][32] = 4'hD;
    SS9[30][32] = 4'hD;
    SS9[31][32] = 4'hE;
    SS9[32][32] = 4'hE;
    SS9[33][32] = 4'hE;
    SS9[34][32] = 4'hE;
    SS9[35][32] = 4'hE;
    SS9[36][32] = 4'hE;
    SS9[37][32] = 4'h0;
    SS9[38][32] = 4'h0;
    SS9[39][32] = 4'h0;
    SS9[40][32] = 4'h0;
    SS9[41][32] = 4'h0;
    SS9[42][32] = 4'h0;
    SS9[43][32] = 4'h0;
    SS9[44][32] = 4'h0;
    SS9[45][32] = 4'h0;
    SS9[46][32] = 4'h0;
    SS9[47][32] = 4'h0;
    SS9[0][33] = 4'h0;
    SS9[1][33] = 4'h0;
    SS9[2][33] = 4'hC;
    SS9[3][33] = 4'hC;
    SS9[4][33] = 4'hC;
    SS9[5][33] = 4'hC;
    SS9[6][33] = 4'hC;
    SS9[7][33] = 4'hC;
    SS9[8][33] = 4'hC;
    SS9[9][33] = 4'hD;
    SS9[10][33] = 4'hD;
    SS9[11][33] = 4'hD;
    SS9[12][33] = 4'hD;
    SS9[13][33] = 4'hD;
    SS9[14][33] = 4'hD;
    SS9[15][33] = 4'hD;
    SS9[16][33] = 4'hD;
    SS9[17][33] = 4'h0;
    SS9[18][33] = 4'h0;
    SS9[19][33] = 4'h0;
    SS9[20][33] = 4'h0;
    SS9[21][33] = 4'hF;
    SS9[22][33] = 4'hD;
    SS9[23][33] = 4'hD;
    SS9[24][33] = 4'h3;
    SS9[25][33] = 4'hD;
    SS9[26][33] = 4'hD;
    SS9[27][33] = 4'hD;
    SS9[28][33] = 4'hD;
    SS9[29][33] = 4'hD;
    SS9[30][33] = 4'hD;
    SS9[31][33] = 4'hE;
    SS9[32][33] = 4'hE;
    SS9[33][33] = 4'hE;
    SS9[34][33] = 4'hE;
    SS9[35][33] = 4'hE;
    SS9[36][33] = 4'hE;
    SS9[37][33] = 4'hE;
    SS9[38][33] = 4'h0;
    SS9[39][33] = 4'h0;
    SS9[40][33] = 4'h0;
    SS9[41][33] = 4'h0;
    SS9[42][33] = 4'h0;
    SS9[43][33] = 4'h0;
    SS9[44][33] = 4'h0;
    SS9[45][33] = 4'h0;
    SS9[46][33] = 4'h0;
    SS9[47][33] = 4'h0;
    SS9[0][34] = 4'h0;
    SS9[1][34] = 4'h0;
    SS9[2][34] = 4'h0;
    SS9[3][34] = 4'hC;
    SS9[4][34] = 4'hC;
    SS9[5][34] = 4'hC;
    SS9[6][34] = 4'h0;
    SS9[7][34] = 4'h0;
    SS9[8][34] = 4'h0;
    SS9[9][34] = 4'hD;
    SS9[10][34] = 4'hD;
    SS9[11][34] = 4'hD;
    SS9[12][34] = 4'hD;
    SS9[13][34] = 4'hD;
    SS9[14][34] = 4'h0;
    SS9[15][34] = 4'h0;
    SS9[16][34] = 4'h0;
    SS9[17][34] = 4'h0;
    SS9[18][34] = 4'h0;
    SS9[19][34] = 4'h0;
    SS9[20][34] = 4'h0;
    SS9[21][34] = 4'h0;
    SS9[22][34] = 4'h3;
    SS9[23][34] = 4'h3;
    SS9[24][34] = 4'h3;
    SS9[25][34] = 4'hD;
    SS9[26][34] = 4'hD;
    SS9[27][34] = 4'hD;
    SS9[28][34] = 4'hD;
    SS9[29][34] = 4'hD;
    SS9[30][34] = 4'hD;
    SS9[31][34] = 4'hD;
    SS9[32][34] = 4'hE;
    SS9[33][34] = 4'hE;
    SS9[34][34] = 4'hE;
    SS9[35][34] = 4'hE;
    SS9[36][34] = 4'hE;
    SS9[37][34] = 4'hE;
    SS9[38][34] = 4'h0;
    SS9[39][34] = 4'h0;
    SS9[40][34] = 4'h0;
    SS9[41][34] = 4'h0;
    SS9[42][34] = 4'h0;
    SS9[43][34] = 4'h0;
    SS9[44][34] = 4'h0;
    SS9[45][34] = 4'h0;
    SS9[46][34] = 4'h0;
    SS9[47][34] = 4'h0;
    SS9[0][35] = 4'h0;
    SS9[1][35] = 4'h0;
    SS9[2][35] = 4'h0;
    SS9[3][35] = 4'hC;
    SS9[4][35] = 4'h0;
    SS9[5][35] = 4'h0;
    SS9[6][35] = 4'h0;
    SS9[7][35] = 4'h0;
    SS9[8][35] = 4'h0;
    SS9[9][35] = 4'hF;
    SS9[10][35] = 4'hD;
    SS9[11][35] = 4'hD;
    SS9[12][35] = 4'h0;
    SS9[13][35] = 4'h0;
    SS9[14][35] = 4'h0;
    SS9[15][35] = 4'h0;
    SS9[16][35] = 4'h0;
    SS9[17][35] = 4'h0;
    SS9[18][35] = 4'h0;
    SS9[19][35] = 4'h0;
    SS9[20][35] = 4'h0;
    SS9[21][35] = 4'h0;
    SS9[22][35] = 4'h3;
    SS9[23][35] = 4'h3;
    SS9[24][35] = 4'h3;
    SS9[25][35] = 4'h3;
    SS9[26][35] = 4'hD;
    SS9[27][35] = 4'h0;
    SS9[28][35] = 4'h0;
    SS9[29][35] = 4'hD;
    SS9[30][35] = 4'hD;
    SS9[31][35] = 4'hD;
    SS9[32][35] = 4'hE;
    SS9[33][35] = 4'hE;
    SS9[34][35] = 4'hE;
    SS9[35][35] = 4'hE;
    SS9[36][35] = 4'hE;
    SS9[37][35] = 4'hE;
    SS9[38][35] = 4'h0;
    SS9[39][35] = 4'h0;
    SS9[40][35] = 4'h0;
    SS9[41][35] = 4'h0;
    SS9[42][35] = 4'h0;
    SS9[43][35] = 4'h0;
    SS9[44][35] = 4'h0;
    SS9[45][35] = 4'h0;
    SS9[46][35] = 4'h0;
    SS9[47][35] = 4'h0;
    SS9[0][36] = 4'h0;
    SS9[1][36] = 4'h0;
    SS9[2][36] = 4'h0;
    SS9[3][36] = 4'h0;
    SS9[4][36] = 4'h0;
    SS9[5][36] = 4'h0;
    SS9[6][36] = 4'h0;
    SS9[7][36] = 4'h0;
    SS9[8][36] = 4'h0;
    SS9[9][36] = 4'h0;
    SS9[10][36] = 4'h0;
    SS9[11][36] = 4'h0;
    SS9[12][36] = 4'h0;
    SS9[13][36] = 4'h0;
    SS9[14][36] = 4'h0;
    SS9[15][36] = 4'h0;
    SS9[16][36] = 4'h0;
    SS9[17][36] = 4'h0;
    SS9[18][36] = 4'h0;
    SS9[19][36] = 4'h0;
    SS9[20][36] = 4'h0;
    SS9[21][36] = 4'h0;
    SS9[22][36] = 4'h0;
    SS9[23][36] = 4'h3;
    SS9[24][36] = 4'h3;
    SS9[25][36] = 4'h0;
    SS9[26][36] = 4'h0;
    SS9[27][36] = 4'h0;
    SS9[28][36] = 4'h0;
    SS9[29][36] = 4'hD;
    SS9[30][36] = 4'hD;
    SS9[31][36] = 4'hD;
    SS9[32][36] = 4'hE;
    SS9[33][36] = 4'hD;
    SS9[34][36] = 4'hD;
    SS9[35][36] = 4'hD;
    SS9[36][36] = 4'hE;
    SS9[37][36] = 4'hE;
    SS9[38][36] = 4'hE;
    SS9[39][36] = 4'h0;
    SS9[40][36] = 4'h0;
    SS9[41][36] = 4'h0;
    SS9[42][36] = 4'h0;
    SS9[43][36] = 4'h0;
    SS9[44][36] = 4'h0;
    SS9[45][36] = 4'h0;
    SS9[46][36] = 4'h0;
    SS9[47][36] = 4'h0;
    SS9[0][37] = 4'h0;
    SS9[1][37] = 4'h0;
    SS9[2][37] = 4'h0;
    SS9[3][37] = 4'h0;
    SS9[4][37] = 4'h0;
    SS9[5][37] = 4'h0;
    SS9[6][37] = 4'h0;
    SS9[7][37] = 4'h0;
    SS9[8][37] = 4'h0;
    SS9[9][37] = 4'h0;
    SS9[10][37] = 4'h0;
    SS9[11][37] = 4'h0;
    SS9[12][37] = 4'h0;
    SS9[13][37] = 4'h0;
    SS9[14][37] = 4'h0;
    SS9[15][37] = 4'h0;
    SS9[16][37] = 4'h0;
    SS9[17][37] = 4'h0;
    SS9[18][37] = 4'h0;
    SS9[19][37] = 4'h0;
    SS9[20][37] = 4'h0;
    SS9[21][37] = 4'h0;
    SS9[22][37] = 4'h0;
    SS9[23][37] = 4'h0;
    SS9[24][37] = 4'h0;
    SS9[25][37] = 4'h0;
    SS9[26][37] = 4'h0;
    SS9[27][37] = 4'h0;
    SS9[28][37] = 4'h0;
    SS9[29][37] = 4'h0;
    SS9[30][37] = 4'h3;
    SS9[31][37] = 4'h3;
    SS9[32][37] = 4'h3;
    SS9[33][37] = 4'hD;
    SS9[34][37] = 4'hD;
    SS9[35][37] = 4'hD;
    SS9[36][37] = 4'hE;
    SS9[37][37] = 4'hE;
    SS9[38][37] = 4'hD;
    SS9[39][37] = 4'h0;
    SS9[40][37] = 4'h0;
    SS9[41][37] = 4'h0;
    SS9[42][37] = 4'h0;
    SS9[43][37] = 4'h0;
    SS9[44][37] = 4'h0;
    SS9[45][37] = 4'h0;
    SS9[46][37] = 4'h0;
    SS9[47][37] = 4'h0;
    SS9[0][38] = 4'h0;
    SS9[1][38] = 4'h0;
    SS9[2][38] = 4'h0;
    SS9[3][38] = 4'h0;
    SS9[4][38] = 4'h0;
    SS9[5][38] = 4'h0;
    SS9[6][38] = 4'h0;
    SS9[7][38] = 4'h0;
    SS9[8][38] = 4'h0;
    SS9[9][38] = 4'h0;
    SS9[10][38] = 4'h0;
    SS9[11][38] = 4'h0;
    SS9[12][38] = 4'h0;
    SS9[13][38] = 4'h0;
    SS9[14][38] = 4'h0;
    SS9[15][38] = 4'h0;
    SS9[16][38] = 4'h0;
    SS9[17][38] = 4'h0;
    SS9[18][38] = 4'h0;
    SS9[19][38] = 4'h0;
    SS9[20][38] = 4'h0;
    SS9[21][38] = 4'h0;
    SS9[22][38] = 4'h0;
    SS9[23][38] = 4'h0;
    SS9[24][38] = 4'h0;
    SS9[25][38] = 4'h0;
    SS9[26][38] = 4'h0;
    SS9[27][38] = 4'h0;
    SS9[28][38] = 4'h0;
    SS9[29][38] = 4'h0;
    SS9[30][38] = 4'h3;
    SS9[31][38] = 4'h3;
    SS9[32][38] = 4'h3;
    SS9[33][38] = 4'hD;
    SS9[34][38] = 4'hD;
    SS9[35][38] = 4'hD;
    SS9[36][38] = 4'hD;
    SS9[37][38] = 4'hD;
    SS9[38][38] = 4'hD;
    SS9[39][38] = 4'hD;
    SS9[40][38] = 4'h0;
    SS9[41][38] = 4'h0;
    SS9[42][38] = 4'h0;
    SS9[43][38] = 4'h0;
    SS9[44][38] = 4'h0;
    SS9[45][38] = 4'h0;
    SS9[46][38] = 4'h0;
    SS9[47][38] = 4'h0;
    SS9[0][39] = 4'h0;
    SS9[1][39] = 4'h0;
    SS9[2][39] = 4'h0;
    SS9[3][39] = 4'h0;
    SS9[4][39] = 4'h0;
    SS9[5][39] = 4'h0;
    SS9[6][39] = 4'h0;
    SS9[7][39] = 4'h0;
    SS9[8][39] = 4'h0;
    SS9[9][39] = 4'h0;
    SS9[10][39] = 4'h0;
    SS9[11][39] = 4'h0;
    SS9[12][39] = 4'h0;
    SS9[13][39] = 4'h0;
    SS9[14][39] = 4'h0;
    SS9[15][39] = 4'h0;
    SS9[16][39] = 4'h0;
    SS9[17][39] = 4'h0;
    SS9[18][39] = 4'h0;
    SS9[19][39] = 4'h0;
    SS9[20][39] = 4'h0;
    SS9[21][39] = 4'h0;
    SS9[22][39] = 4'h0;
    SS9[23][39] = 4'h0;
    SS9[24][39] = 4'h0;
    SS9[25][39] = 4'h0;
    SS9[26][39] = 4'h0;
    SS9[27][39] = 4'h0;
    SS9[28][39] = 4'h0;
    SS9[29][39] = 4'h0;
    SS9[30][39] = 4'h3;
    SS9[31][39] = 4'h3;
    SS9[32][39] = 4'h3;
    SS9[33][39] = 4'h0;
    SS9[34][39] = 4'hD;
    SS9[35][39] = 4'hD;
    SS9[36][39] = 4'hD;
    SS9[37][39] = 4'hD;
    SS9[38][39] = 4'hD;
    SS9[39][39] = 4'hD;
    SS9[40][39] = 4'h0;
    SS9[41][39] = 4'h0;
    SS9[42][39] = 4'h0;
    SS9[43][39] = 4'h0;
    SS9[44][39] = 4'h0;
    SS9[45][39] = 4'h0;
    SS9[46][39] = 4'h0;
    SS9[47][39] = 4'h0;
    SS9[0][40] = 4'h0;
    SS9[1][40] = 4'h0;
    SS9[2][40] = 4'h0;
    SS9[3][40] = 4'h0;
    SS9[4][40] = 4'h0;
    SS9[5][40] = 4'h0;
    SS9[6][40] = 4'h0;
    SS9[7][40] = 4'h0;
    SS9[8][40] = 4'h0;
    SS9[9][40] = 4'h0;
    SS9[10][40] = 4'h0;
    SS9[11][40] = 4'h0;
    SS9[12][40] = 4'h0;
    SS9[13][40] = 4'h0;
    SS9[14][40] = 4'h0;
    SS9[15][40] = 4'h0;
    SS9[16][40] = 4'h0;
    SS9[17][40] = 4'h0;
    SS9[18][40] = 4'h0;
    SS9[19][40] = 4'h0;
    SS9[20][40] = 4'h0;
    SS9[21][40] = 4'h0;
    SS9[22][40] = 4'h0;
    SS9[23][40] = 4'h0;
    SS9[24][40] = 4'h0;
    SS9[25][40] = 4'h0;
    SS9[26][40] = 4'h0;
    SS9[27][40] = 4'h0;
    SS9[28][40] = 4'h0;
    SS9[29][40] = 4'h0;
    SS9[30][40] = 4'h0;
    SS9[31][40] = 4'h0;
    SS9[32][40] = 4'h0;
    SS9[33][40] = 4'h0;
    SS9[34][40] = 4'hD;
    SS9[35][40] = 4'hD;
    SS9[36][40] = 4'hD;
    SS9[37][40] = 4'hD;
    SS9[38][40] = 4'hD;
    SS9[39][40] = 4'hD;
    SS9[40][40] = 4'h0;
    SS9[41][40] = 4'h0;
    SS9[42][40] = 4'h0;
    SS9[43][40] = 4'h0;
    SS9[44][40] = 4'h0;
    SS9[45][40] = 4'h0;
    SS9[46][40] = 4'h0;
    SS9[47][40] = 4'h0;
    SS9[0][41] = 4'h0;
    SS9[1][41] = 4'h0;
    SS9[2][41] = 4'h0;
    SS9[3][41] = 4'h0;
    SS9[4][41] = 4'h0;
    SS9[5][41] = 4'h0;
    SS9[6][41] = 4'h0;
    SS9[7][41] = 4'h0;
    SS9[8][41] = 4'h0;
    SS9[9][41] = 4'h0;
    SS9[10][41] = 4'h0;
    SS9[11][41] = 4'h0;
    SS9[12][41] = 4'h0;
    SS9[13][41] = 4'h0;
    SS9[14][41] = 4'h0;
    SS9[15][41] = 4'h0;
    SS9[16][41] = 4'h0;
    SS9[17][41] = 4'h0;
    SS9[18][41] = 4'h0;
    SS9[19][41] = 4'h0;
    SS9[20][41] = 4'h0;
    SS9[21][41] = 4'h0;
    SS9[22][41] = 4'h0;
    SS9[23][41] = 4'h0;
    SS9[24][41] = 4'h0;
    SS9[25][41] = 4'h0;
    SS9[26][41] = 4'h0;
    SS9[27][41] = 4'h0;
    SS9[28][41] = 4'h0;
    SS9[29][41] = 4'h0;
    SS9[30][41] = 4'h0;
    SS9[31][41] = 4'h0;
    SS9[32][41] = 4'h0;
    SS9[33][41] = 4'h0;
    SS9[34][41] = 4'hD;
    SS9[35][41] = 4'hD;
    SS9[36][41] = 4'h0;
    SS9[37][41] = 4'h0;
    SS9[38][41] = 4'hD;
    SS9[39][41] = 4'hD;
    SS9[40][41] = 4'hD;
    SS9[41][41] = 4'h0;
    SS9[42][41] = 4'h0;
    SS9[43][41] = 4'h0;
    SS9[44][41] = 4'h0;
    SS9[45][41] = 4'h0;
    SS9[46][41] = 4'h0;
    SS9[47][41] = 4'h0;
    SS9[0][42] = 4'h0;
    SS9[1][42] = 4'h0;
    SS9[2][42] = 4'h0;
    SS9[3][42] = 4'h0;
    SS9[4][42] = 4'h0;
    SS9[5][42] = 4'h0;
    SS9[6][42] = 4'h0;
    SS9[7][42] = 4'h0;
    SS9[8][42] = 4'h0;
    SS9[9][42] = 4'h0;
    SS9[10][42] = 4'h0;
    SS9[11][42] = 4'h0;
    SS9[12][42] = 4'h0;
    SS9[13][42] = 4'h0;
    SS9[14][42] = 4'h0;
    SS9[15][42] = 4'h0;
    SS9[16][42] = 4'h0;
    SS9[17][42] = 4'h0;
    SS9[18][42] = 4'h0;
    SS9[19][42] = 4'h0;
    SS9[20][42] = 4'h0;
    SS9[21][42] = 4'h0;
    SS9[22][42] = 4'h0;
    SS9[23][42] = 4'h0;
    SS9[24][42] = 4'h0;
    SS9[25][42] = 4'h0;
    SS9[26][42] = 4'h0;
    SS9[27][42] = 4'h0;
    SS9[28][42] = 4'h0;
    SS9[29][42] = 4'h0;
    SS9[30][42] = 4'h0;
    SS9[31][42] = 4'h0;
    SS9[32][42] = 4'h0;
    SS9[33][42] = 4'h0;
    SS9[34][42] = 4'h0;
    SS9[35][42] = 4'h0;
    SS9[36][42] = 4'h0;
    SS9[37][42] = 4'h0;
    SS9[38][42] = 4'hD;
    SS9[39][42] = 4'hD;
    SS9[40][42] = 4'hD;
    SS9[41][42] = 4'h0;
    SS9[42][42] = 4'h0;
    SS9[43][42] = 4'h0;
    SS9[44][42] = 4'h0;
    SS9[45][42] = 4'h0;
    SS9[46][42] = 4'h0;
    SS9[47][42] = 4'h0;
    SS9[0][43] = 4'h0;
    SS9[1][43] = 4'h0;
    SS9[2][43] = 4'h0;
    SS9[3][43] = 4'h0;
    SS9[4][43] = 4'h0;
    SS9[5][43] = 4'h0;
    SS9[6][43] = 4'h0;
    SS9[7][43] = 4'h0;
    SS9[8][43] = 4'h0;
    SS9[9][43] = 4'h0;
    SS9[10][43] = 4'h0;
    SS9[11][43] = 4'h0;
    SS9[12][43] = 4'h0;
    SS9[13][43] = 4'h0;
    SS9[14][43] = 4'h0;
    SS9[15][43] = 4'h0;
    SS9[16][43] = 4'h0;
    SS9[17][43] = 4'h0;
    SS9[18][43] = 4'h0;
    SS9[19][43] = 4'h0;
    SS9[20][43] = 4'h0;
    SS9[21][43] = 4'h0;
    SS9[22][43] = 4'h0;
    SS9[23][43] = 4'h0;
    SS9[24][43] = 4'h0;
    SS9[25][43] = 4'h0;
    SS9[26][43] = 4'h0;
    SS9[27][43] = 4'h0;
    SS9[28][43] = 4'h0;
    SS9[29][43] = 4'h0;
    SS9[30][43] = 4'h0;
    SS9[31][43] = 4'h0;
    SS9[32][43] = 4'h0;
    SS9[33][43] = 4'h0;
    SS9[34][43] = 4'h0;
    SS9[35][43] = 4'h0;
    SS9[36][43] = 4'h0;
    SS9[37][43] = 4'h0;
    SS9[38][43] = 4'hD;
    SS9[39][43] = 4'h0;
    SS9[40][43] = 4'h0;
    SS9[41][43] = 4'h0;
    SS9[42][43] = 4'h0;
    SS9[43][43] = 4'h0;
    SS9[44][43] = 4'h0;
    SS9[45][43] = 4'h0;
    SS9[46][43] = 4'h0;
    SS9[47][43] = 4'h0;
    SS9[0][44] = 4'h0;
    SS9[1][44] = 4'h0;
    SS9[2][44] = 4'h0;
    SS9[3][44] = 4'h0;
    SS9[4][44] = 4'h0;
    SS9[5][44] = 4'h0;
    SS9[6][44] = 4'h0;
    SS9[7][44] = 4'h0;
    SS9[8][44] = 4'h0;
    SS9[9][44] = 4'h0;
    SS9[10][44] = 4'h0;
    SS9[11][44] = 4'h0;
    SS9[12][44] = 4'h0;
    SS9[13][44] = 4'h0;
    SS9[14][44] = 4'h0;
    SS9[15][44] = 4'h0;
    SS9[16][44] = 4'h0;
    SS9[17][44] = 4'h0;
    SS9[18][44] = 4'h0;
    SS9[19][44] = 4'h0;
    SS9[20][44] = 4'h0;
    SS9[21][44] = 4'h0;
    SS9[22][44] = 4'h0;
    SS9[23][44] = 4'h0;
    SS9[24][44] = 4'h0;
    SS9[25][44] = 4'h0;
    SS9[26][44] = 4'h0;
    SS9[27][44] = 4'h0;
    SS9[28][44] = 4'h0;
    SS9[29][44] = 4'h0;
    SS9[30][44] = 4'h0;
    SS9[31][44] = 4'h0;
    SS9[32][44] = 4'h0;
    SS9[33][44] = 4'h0;
    SS9[34][44] = 4'h0;
    SS9[35][44] = 4'h0;
    SS9[36][44] = 4'h0;
    SS9[37][44] = 4'h0;
    SS9[38][44] = 4'h0;
    SS9[39][44] = 4'h0;
    SS9[40][44] = 4'h0;
    SS9[41][44] = 4'h0;
    SS9[42][44] = 4'h0;
    SS9[43][44] = 4'h0;
    SS9[44][44] = 4'h0;
    SS9[45][44] = 4'h0;
    SS9[46][44] = 4'h0;
    SS9[47][44] = 4'h0;
    SS9[0][45] = 4'h0;
    SS9[1][45] = 4'h0;
    SS9[2][45] = 4'h0;
    SS9[3][45] = 4'h0;
    SS9[4][45] = 4'h0;
    SS9[5][45] = 4'h0;
    SS9[6][45] = 4'h0;
    SS9[7][45] = 4'h0;
    SS9[8][45] = 4'h0;
    SS9[9][45] = 4'h0;
    SS9[10][45] = 4'h0;
    SS9[11][45] = 4'h0;
    SS9[12][45] = 4'h0;
    SS9[13][45] = 4'h0;
    SS9[14][45] = 4'h0;
    SS9[15][45] = 4'h0;
    SS9[16][45] = 4'h0;
    SS9[17][45] = 4'h0;
    SS9[18][45] = 4'h0;
    SS9[19][45] = 4'h0;
    SS9[20][45] = 4'h0;
    SS9[21][45] = 4'h0;
    SS9[22][45] = 4'h0;
    SS9[23][45] = 4'h0;
    SS9[24][45] = 4'h0;
    SS9[25][45] = 4'h0;
    SS9[26][45] = 4'h0;
    SS9[27][45] = 4'h0;
    SS9[28][45] = 4'h0;
    SS9[29][45] = 4'h0;
    SS9[30][45] = 4'h0;
    SS9[31][45] = 4'h0;
    SS9[32][45] = 4'h0;
    SS9[33][45] = 4'h0;
    SS9[34][45] = 4'h0;
    SS9[35][45] = 4'h0;
    SS9[36][45] = 4'h0;
    SS9[37][45] = 4'h0;
    SS9[38][45] = 4'h0;
    SS9[39][45] = 4'h0;
    SS9[40][45] = 4'h0;
    SS9[41][45] = 4'h0;
    SS9[42][45] = 4'h0;
    SS9[43][45] = 4'h0;
    SS9[44][45] = 4'h0;
    SS9[45][45] = 4'h0;
    SS9[46][45] = 4'h0;
    SS9[47][45] = 4'h0;
    SS9[0][46] = 4'h0;
    SS9[1][46] = 4'h0;
    SS9[2][46] = 4'h0;
    SS9[3][46] = 4'h0;
    SS9[4][46] = 4'h0;
    SS9[5][46] = 4'h0;
    SS9[6][46] = 4'h0;
    SS9[7][46] = 4'h0;
    SS9[8][46] = 4'h0;
    SS9[9][46] = 4'h0;
    SS9[10][46] = 4'h0;
    SS9[11][46] = 4'h0;
    SS9[12][46] = 4'h0;
    SS9[13][46] = 4'h0;
    SS9[14][46] = 4'h0;
    SS9[15][46] = 4'h0;
    SS9[16][46] = 4'h0;
    SS9[17][46] = 4'h0;
    SS9[18][46] = 4'h0;
    SS9[19][46] = 4'h0;
    SS9[20][46] = 4'h0;
    SS9[21][46] = 4'h0;
    SS9[22][46] = 4'h0;
    SS9[23][46] = 4'h0;
    SS9[24][46] = 4'h0;
    SS9[25][46] = 4'h0;
    SS9[26][46] = 4'h0;
    SS9[27][46] = 4'h0;
    SS9[28][46] = 4'h0;
    SS9[29][46] = 4'h0;
    SS9[30][46] = 4'h0;
    SS9[31][46] = 4'h0;
    SS9[32][46] = 4'h0;
    SS9[33][46] = 4'h0;
    SS9[34][46] = 4'h0;
    SS9[35][46] = 4'h0;
    SS9[36][46] = 4'h0;
    SS9[37][46] = 4'h0;
    SS9[38][46] = 4'h0;
    SS9[39][46] = 4'h0;
    SS9[40][46] = 4'h0;
    SS9[41][46] = 4'h0;
    SS9[42][46] = 4'h0;
    SS9[43][46] = 4'h0;
    SS9[44][46] = 4'h0;
    SS9[45][46] = 4'h0;
    SS9[46][46] = 4'h0;
    SS9[47][46] = 4'h0;
    SS9[0][47] = 4'h0;
    SS9[1][47] = 4'h0;
    SS9[2][47] = 4'h0;
    SS9[3][47] = 4'h0;
    SS9[4][47] = 4'h0;
    SS9[5][47] = 4'h0;
    SS9[6][47] = 4'h0;
    SS9[7][47] = 4'h0;
    SS9[8][47] = 4'h0;
    SS9[9][47] = 4'h0;
    SS9[10][47] = 4'h0;
    SS9[11][47] = 4'h0;
    SS9[12][47] = 4'h0;
    SS9[13][47] = 4'h0;
    SS9[14][47] = 4'h0;
    SS9[15][47] = 4'h0;
    SS9[16][47] = 4'h0;
    SS9[17][47] = 4'h0;
    SS9[18][47] = 4'h0;
    SS9[19][47] = 4'h0;
    SS9[20][47] = 4'h0;
    SS9[21][47] = 4'h0;
    SS9[22][47] = 4'h0;
    SS9[23][47] = 4'h0;
    SS9[24][47] = 4'h0;
    SS9[25][47] = 4'h0;
    SS9[26][47] = 4'h0;
    SS9[27][47] = 4'h0;
    SS9[28][47] = 4'h0;
    SS9[29][47] = 4'h0;
    SS9[30][47] = 4'h0;
    SS9[31][47] = 4'h0;
    SS9[32][47] = 4'h0;
    SS9[33][47] = 4'h0;
    SS9[34][47] = 4'h0;
    SS9[35][47] = 4'h0;
    SS9[36][47] = 4'h0;
    SS9[37][47] = 4'h0;
    SS9[38][47] = 4'h0;
    SS9[39][47] = 4'h0;
    SS9[40][47] = 4'h0;
    SS9[41][47] = 4'h0;
    SS9[42][47] = 4'h0;
    SS9[43][47] = 4'h0;
    SS9[44][47] = 4'h0;
    SS9[45][47] = 4'h0;
    SS9[46][47] = 4'h0;
    SS9[47][47] = 4'h0;
 
//SS 10
    SS10[0][0] = 4'h0;
    SS10[1][0] = 4'h0;
    SS10[2][0] = 4'h0;
    SS10[3][0] = 4'h0;
    SS10[4][0] = 4'h0;
    SS10[5][0] = 4'h0;
    SS10[6][0] = 4'h0;
    SS10[7][0] = 4'h0;
    SS10[8][0] = 4'h0;
    SS10[9][0] = 4'h0;
    SS10[10][0] = 4'h0;
    SS10[11][0] = 4'h0;
    SS10[12][0] = 4'h0;
    SS10[13][0] = 4'h0;
    SS10[14][0] = 4'h0;
    SS10[15][0] = 4'h0;
    SS10[16][0] = 4'h0;
    SS10[17][0] = 4'h0;
    SS10[18][0] = 4'h0;
    SS10[19][0] = 4'h0;
    SS10[20][0] = 4'h0;
    SS10[21][0] = 4'h0;
    SS10[22][0] = 4'h0;
    SS10[23][0] = 4'h0;
    SS10[24][0] = 4'h0;
    SS10[25][0] = 4'h0;
    SS10[26][0] = 4'h0;
    SS10[27][0] = 4'h0;
    SS10[28][0] = 4'h0;
    SS10[29][0] = 4'h0;
    SS10[30][0] = 4'hD;
    SS10[31][0] = 4'hD;
    SS10[32][0] = 4'hD;
    SS10[33][0] = 4'h0;
    SS10[34][0] = 4'h0;
    SS10[35][0] = 4'h0;
    SS10[36][0] = 4'h0;
    SS10[37][0] = 4'h0;
    SS10[38][0] = 4'h0;
    SS10[39][0] = 4'h0;
    SS10[40][0] = 4'h0;
    SS10[41][0] = 4'h0;
    SS10[42][0] = 4'h0;
    SS10[43][0] = 4'h0;
    SS10[44][0] = 4'h0;
    SS10[45][0] = 4'h0;
    SS10[46][0] = 4'h0;
    SS10[47][0] = 4'h0;
    SS10[0][1] = 4'h0;
    SS10[1][1] = 4'h0;
    SS10[2][1] = 4'h0;
    SS10[3][1] = 4'h0;
    SS10[4][1] = 4'h0;
    SS10[5][1] = 4'h0;
    SS10[6][1] = 4'h0;
    SS10[7][1] = 4'h0;
    SS10[8][1] = 4'h0;
    SS10[9][1] = 4'h0;
    SS10[10][1] = 4'h0;
    SS10[11][1] = 4'h0;
    SS10[12][1] = 4'h0;
    SS10[13][1] = 4'h0;
    SS10[14][1] = 4'h0;
    SS10[15][1] = 4'h0;
    SS10[16][1] = 4'h0;
    SS10[17][1] = 4'h0;
    SS10[18][1] = 4'h0;
    SS10[19][1] = 4'h0;
    SS10[20][1] = 4'h0;
    SS10[21][1] = 4'h0;
    SS10[22][1] = 4'h0;
    SS10[23][1] = 4'h0;
    SS10[24][1] = 4'h0;
    SS10[25][1] = 4'h0;
    SS10[26][1] = 4'h0;
    SS10[27][1] = 4'h0;
    SS10[28][1] = 4'h0;
    SS10[29][1] = 4'h0;
    SS10[30][1] = 4'hD;
    SS10[31][1] = 4'hD;
    SS10[32][1] = 4'hD;
    SS10[33][1] = 4'h0;
    SS10[34][1] = 4'h0;
    SS10[35][1] = 4'h0;
    SS10[36][1] = 4'h0;
    SS10[37][1] = 4'h0;
    SS10[38][1] = 4'h0;
    SS10[39][1] = 4'h0;
    SS10[40][1] = 4'h0;
    SS10[41][1] = 4'h0;
    SS10[42][1] = 4'h0;
    SS10[43][1] = 4'h0;
    SS10[44][1] = 4'h0;
    SS10[45][1] = 4'h0;
    SS10[46][1] = 4'h0;
    SS10[47][1] = 4'h0;
    SS10[0][2] = 4'h0;
    SS10[1][2] = 4'h0;
    SS10[2][2] = 4'h0;
    SS10[3][2] = 4'h0;
    SS10[4][2] = 4'h0;
    SS10[5][2] = 4'h0;
    SS10[6][2] = 4'h0;
    SS10[7][2] = 4'h0;
    SS10[8][2] = 4'h0;
    SS10[9][2] = 4'h0;
    SS10[10][2] = 4'h0;
    SS10[11][2] = 4'h0;
    SS10[12][2] = 4'h0;
    SS10[13][2] = 4'h0;
    SS10[14][2] = 4'h0;
    SS10[15][2] = 4'h0;
    SS10[16][2] = 4'h0;
    SS10[17][2] = 4'h0;
    SS10[18][2] = 4'h0;
    SS10[19][2] = 4'h0;
    SS10[20][2] = 4'h0;
    SS10[21][2] = 4'h0;
    SS10[22][2] = 4'h0;
    SS10[23][2] = 4'h0;
    SS10[24][2] = 4'h0;
    SS10[25][2] = 4'h0;
    SS10[26][2] = 4'h0;
    SS10[27][2] = 4'h0;
    SS10[28][2] = 4'h0;
    SS10[29][2] = 4'h0;
    SS10[30][2] = 4'hD;
    SS10[31][2] = 4'hD;
    SS10[32][2] = 4'hD;
    SS10[33][2] = 4'h0;
    SS10[34][2] = 4'h0;
    SS10[35][2] = 4'h0;
    SS10[36][2] = 4'h0;
    SS10[37][2] = 4'h0;
    SS10[38][2] = 4'h0;
    SS10[39][2] = 4'h0;
    SS10[40][2] = 4'h0;
    SS10[41][2] = 4'h0;
    SS10[42][2] = 4'h0;
    SS10[43][2] = 4'h0;
    SS10[44][2] = 4'h0;
    SS10[45][2] = 4'h0;
    SS10[46][2] = 4'h0;
    SS10[47][2] = 4'h0;
    SS10[0][3] = 4'h0;
    SS10[1][3] = 4'h0;
    SS10[2][3] = 4'h0;
    SS10[3][3] = 4'h0;
    SS10[4][3] = 4'h0;
    SS10[5][3] = 4'h0;
    SS10[6][3] = 4'h0;
    SS10[7][3] = 4'h0;
    SS10[8][3] = 4'h0;
    SS10[9][3] = 4'h0;
    SS10[10][3] = 4'h0;
    SS10[11][3] = 4'h0;
    SS10[12][3] = 4'h0;
    SS10[13][3] = 4'h0;
    SS10[14][3] = 4'h0;
    SS10[15][3] = 4'h0;
    SS10[16][3] = 4'h0;
    SS10[17][3] = 4'h0;
    SS10[18][3] = 4'h0;
    SS10[19][3] = 4'h0;
    SS10[20][3] = 4'h0;
    SS10[21][3] = 4'h0;
    SS10[22][3] = 4'h0;
    SS10[23][3] = 4'h0;
    SS10[24][3] = 4'h0;
    SS10[25][3] = 4'h0;
    SS10[26][3] = 4'h0;
    SS10[27][3] = 4'hD;
    SS10[28][3] = 4'hD;
    SS10[29][3] = 4'hD;
    SS10[30][3] = 4'hD;
    SS10[31][3] = 4'hD;
    SS10[32][3] = 4'hD;
    SS10[33][3] = 4'h0;
    SS10[34][3] = 4'h0;
    SS10[35][3] = 4'h0;
    SS10[36][3] = 4'h0;
    SS10[37][3] = 4'h0;
    SS10[38][3] = 4'h0;
    SS10[39][3] = 4'h0;
    SS10[40][3] = 4'h0;
    SS10[41][3] = 4'h0;
    SS10[42][3] = 4'h0;
    SS10[43][3] = 4'h0;
    SS10[44][3] = 4'h0;
    SS10[45][3] = 4'h0;
    SS10[46][3] = 4'h0;
    SS10[47][3] = 4'h0;
    SS10[0][4] = 4'h0;
    SS10[1][4] = 4'h0;
    SS10[2][4] = 4'h0;
    SS10[3][4] = 4'h0;
    SS10[4][4] = 4'h0;
    SS10[5][4] = 4'h0;
    SS10[6][4] = 4'h0;
    SS10[7][4] = 4'h0;
    SS10[8][4] = 4'h0;
    SS10[9][4] = 4'h0;
    SS10[10][4] = 4'h0;
    SS10[11][4] = 4'h0;
    SS10[12][4] = 4'h0;
    SS10[13][4] = 4'h0;
    SS10[14][4] = 4'h0;
    SS10[15][4] = 4'h0;
    SS10[16][4] = 4'h0;
    SS10[17][4] = 4'h0;
    SS10[18][4] = 4'h0;
    SS10[19][4] = 4'h0;
    SS10[20][4] = 4'h0;
    SS10[21][4] = 4'h0;
    SS10[22][4] = 4'h0;
    SS10[23][4] = 4'h0;
    SS10[24][4] = 4'h0;
    SS10[25][4] = 4'h0;
    SS10[26][4] = 4'h0;
    SS10[27][4] = 4'hD;
    SS10[28][4] = 4'hD;
    SS10[29][4] = 4'hD;
    SS10[30][4] = 4'hD;
    SS10[31][4] = 4'hD;
    SS10[32][4] = 4'hD;
    SS10[33][4] = 4'h0;
    SS10[34][4] = 4'h0;
    SS10[35][4] = 4'h0;
    SS10[36][4] = 4'h0;
    SS10[37][4] = 4'h0;
    SS10[38][4] = 4'h0;
    SS10[39][4] = 4'h0;
    SS10[40][4] = 4'h0;
    SS10[41][4] = 4'h0;
    SS10[42][4] = 4'h0;
    SS10[43][4] = 4'h0;
    SS10[44][4] = 4'h0;
    SS10[45][4] = 4'h0;
    SS10[46][4] = 4'h0;
    SS10[47][4] = 4'h0;
    SS10[0][5] = 4'h0;
    SS10[1][5] = 4'h0;
    SS10[2][5] = 4'h0;
    SS10[3][5] = 4'h0;
    SS10[4][5] = 4'h0;
    SS10[5][5] = 4'h0;
    SS10[6][5] = 4'h0;
    SS10[7][5] = 4'h0;
    SS10[8][5] = 4'h0;
    SS10[9][5] = 4'h0;
    SS10[10][5] = 4'h0;
    SS10[11][5] = 4'h0;
    SS10[12][5] = 4'h0;
    SS10[13][5] = 4'h0;
    SS10[14][5] = 4'h0;
    SS10[15][5] = 4'h0;
    SS10[16][5] = 4'h0;
    SS10[17][5] = 4'h0;
    SS10[18][5] = 4'h0;
    SS10[19][5] = 4'h0;
    SS10[20][5] = 4'h0;
    SS10[21][5] = 4'h0;
    SS10[22][5] = 4'h0;
    SS10[23][5] = 4'h0;
    SS10[24][5] = 4'h0;
    SS10[25][5] = 4'h0;
    SS10[26][5] = 4'h0;
    SS10[27][5] = 4'hD;
    SS10[28][5] = 4'hD;
    SS10[29][5] = 4'hD;
    SS10[30][5] = 4'hD;
    SS10[31][5] = 4'hD;
    SS10[32][5] = 4'hD;
    SS10[33][5] = 4'h0;
    SS10[34][5] = 4'h0;
    SS10[35][5] = 4'h0;
    SS10[36][5] = 4'h0;
    SS10[37][5] = 4'h0;
    SS10[38][5] = 4'h0;
    SS10[39][5] = 4'h0;
    SS10[40][5] = 4'h0;
    SS10[41][5] = 4'h0;
    SS10[42][5] = 4'h0;
    SS10[43][5] = 4'h0;
    SS10[44][5] = 4'h0;
    SS10[45][5] = 4'h0;
    SS10[46][5] = 4'h0;
    SS10[47][5] = 4'h0;
    SS10[0][6] = 4'h0;
    SS10[1][6] = 4'h0;
    SS10[2][6] = 4'h0;
    SS10[3][6] = 4'h0;
    SS10[4][6] = 4'h0;
    SS10[5][6] = 4'h0;
    SS10[6][6] = 4'h0;
    SS10[7][6] = 4'h0;
    SS10[8][6] = 4'h0;
    SS10[9][6] = 4'h0;
    SS10[10][6] = 4'h0;
    SS10[11][6] = 4'h0;
    SS10[12][6] = 4'h0;
    SS10[13][6] = 4'h0;
    SS10[14][6] = 4'h0;
    SS10[15][6] = 4'h0;
    SS10[16][6] = 4'h0;
    SS10[17][6] = 4'h0;
    SS10[18][6] = 4'h0;
    SS10[19][6] = 4'h0;
    SS10[20][6] = 4'h0;
    SS10[21][6] = 4'h0;
    SS10[22][6] = 4'h0;
    SS10[23][6] = 4'h0;
    SS10[24][6] = 4'h3;
    SS10[25][6] = 4'h3;
    SS10[26][6] = 4'h3;
    SS10[27][6] = 4'hD;
    SS10[28][6] = 4'hD;
    SS10[29][6] = 4'hD;
    SS10[30][6] = 4'hE;
    SS10[31][6] = 4'hE;
    SS10[32][6] = 4'hE;
    SS10[33][6] = 4'h0;
    SS10[34][6] = 4'h0;
    SS10[35][6] = 4'h0;
    SS10[36][6] = 4'h0;
    SS10[37][6] = 4'h0;
    SS10[38][6] = 4'h0;
    SS10[39][6] = 4'h0;
    SS10[40][6] = 4'h0;
    SS10[41][6] = 4'h0;
    SS10[42][6] = 4'h0;
    SS10[43][6] = 4'h0;
    SS10[44][6] = 4'h0;
    SS10[45][6] = 4'h0;
    SS10[46][6] = 4'h0;
    SS10[47][6] = 4'h0;
    SS10[0][7] = 4'h0;
    SS10[1][7] = 4'h0;
    SS10[2][7] = 4'h0;
    SS10[3][7] = 4'h0;
    SS10[4][7] = 4'h0;
    SS10[5][7] = 4'h0;
    SS10[6][7] = 4'h0;
    SS10[7][7] = 4'h0;
    SS10[8][7] = 4'h0;
    SS10[9][7] = 4'h0;
    SS10[10][7] = 4'h0;
    SS10[11][7] = 4'h0;
    SS10[12][7] = 4'h0;
    SS10[13][7] = 4'h0;
    SS10[14][7] = 4'h0;
    SS10[15][7] = 4'h0;
    SS10[16][7] = 4'h0;
    SS10[17][7] = 4'h0;
    SS10[18][7] = 4'h0;
    SS10[19][7] = 4'h0;
    SS10[20][7] = 4'h0;
    SS10[21][7] = 4'h0;
    SS10[22][7] = 4'h0;
    SS10[23][7] = 4'h0;
    SS10[24][7] = 4'h3;
    SS10[25][7] = 4'h3;
    SS10[26][7] = 4'h3;
    SS10[27][7] = 4'hD;
    SS10[28][7] = 4'hD;
    SS10[29][7] = 4'hD;
    SS10[30][7] = 4'hE;
    SS10[31][7] = 4'hE;
    SS10[32][7] = 4'hE;
    SS10[33][7] = 4'h0;
    SS10[34][7] = 4'h0;
    SS10[35][7] = 4'h0;
    SS10[36][7] = 4'h0;
    SS10[37][7] = 4'h0;
    SS10[38][7] = 4'h0;
    SS10[39][7] = 4'h0;
    SS10[40][7] = 4'h0;
    SS10[41][7] = 4'h0;
    SS10[42][7] = 4'h0;
    SS10[43][7] = 4'h0;
    SS10[44][7] = 4'h0;
    SS10[45][7] = 4'h0;
    SS10[46][7] = 4'h0;
    SS10[47][7] = 4'h0;
    SS10[0][8] = 4'h0;
    SS10[1][8] = 4'h0;
    SS10[2][8] = 4'h0;
    SS10[3][8] = 4'h0;
    SS10[4][8] = 4'h0;
    SS10[5][8] = 4'h0;
    SS10[6][8] = 4'h0;
    SS10[7][8] = 4'h0;
    SS10[8][8] = 4'h0;
    SS10[9][8] = 4'h0;
    SS10[10][8] = 4'h0;
    SS10[11][8] = 4'h0;
    SS10[12][8] = 4'h0;
    SS10[13][8] = 4'h0;
    SS10[14][8] = 4'h0;
    SS10[15][8] = 4'h0;
    SS10[16][8] = 4'h0;
    SS10[17][8] = 4'h0;
    SS10[18][8] = 4'h0;
    SS10[19][8] = 4'h0;
    SS10[20][8] = 4'h0;
    SS10[21][8] = 4'h0;
    SS10[22][8] = 4'h0;
    SS10[23][8] = 4'h0;
    SS10[24][8] = 4'h3;
    SS10[25][8] = 4'h3;
    SS10[26][8] = 4'h3;
    SS10[27][8] = 4'hD;
    SS10[28][8] = 4'hD;
    SS10[29][8] = 4'hD;
    SS10[30][8] = 4'hE;
    SS10[31][8] = 4'hE;
    SS10[32][8] = 4'hE;
    SS10[33][8] = 4'h0;
    SS10[34][8] = 4'h0;
    SS10[35][8] = 4'h0;
    SS10[36][8] = 4'h0;
    SS10[37][8] = 4'h0;
    SS10[38][8] = 4'h0;
    SS10[39][8] = 4'h0;
    SS10[40][8] = 4'h0;
    SS10[41][8] = 4'h0;
    SS10[42][8] = 4'h0;
    SS10[43][8] = 4'h0;
    SS10[44][8] = 4'h0;
    SS10[45][8] = 4'h0;
    SS10[46][8] = 4'h0;
    SS10[47][8] = 4'h0;
    SS10[0][9] = 4'h0;
    SS10[1][9] = 4'h0;
    SS10[2][9] = 4'h0;
    SS10[3][9] = 4'h0;
    SS10[4][9] = 4'h0;
    SS10[5][9] = 4'h0;
    SS10[6][9] = 4'h0;
    SS10[7][9] = 4'h0;
    SS10[8][9] = 4'h0;
    SS10[9][9] = 4'h0;
    SS10[10][9] = 4'h0;
    SS10[11][9] = 4'h0;
    SS10[12][9] = 4'h0;
    SS10[13][9] = 4'h0;
    SS10[14][9] = 4'h0;
    SS10[15][9] = 4'h0;
    SS10[16][9] = 4'h0;
    SS10[17][9] = 4'h0;
    SS10[18][9] = 4'h0;
    SS10[19][9] = 4'h0;
    SS10[20][9] = 4'h0;
    SS10[21][9] = 4'h0;
    SS10[22][9] = 4'h0;
    SS10[23][9] = 4'h0;
    SS10[24][9] = 4'hD;
    SS10[25][9] = 4'hD;
    SS10[26][9] = 4'hD;
    SS10[27][9] = 4'hE;
    SS10[28][9] = 4'hE;
    SS10[29][9] = 4'hE;
    SS10[30][9] = 4'hE;
    SS10[31][9] = 4'hE;
    SS10[32][9] = 4'hE;
    SS10[33][9] = 4'h0;
    SS10[34][9] = 4'h0;
    SS10[35][9] = 4'h0;
    SS10[36][9] = 4'h0;
    SS10[37][9] = 4'h0;
    SS10[38][9] = 4'h0;
    SS10[39][9] = 4'hC;
    SS10[40][9] = 4'hC;
    SS10[41][9] = 4'hC;
    SS10[42][9] = 4'hC;
    SS10[43][9] = 4'hC;
    SS10[44][9] = 4'hC;
    SS10[45][9] = 4'hD;
    SS10[46][9] = 4'hD;
    SS10[47][9] = 4'hD;
    SS10[0][10] = 4'h0;
    SS10[1][10] = 4'h0;
    SS10[2][10] = 4'h0;
    SS10[3][10] = 4'h0;
    SS10[4][10] = 4'h0;
    SS10[5][10] = 4'h0;
    SS10[6][10] = 4'h0;
    SS10[7][10] = 4'h0;
    SS10[8][10] = 4'h0;
    SS10[9][10] = 4'h0;
    SS10[10][10] = 4'h0;
    SS10[11][10] = 4'h0;
    SS10[12][10] = 4'h0;
    SS10[13][10] = 4'h0;
    SS10[14][10] = 4'h0;
    SS10[15][10] = 4'h0;
    SS10[16][10] = 4'h0;
    SS10[17][10] = 4'h0;
    SS10[18][10] = 4'h0;
    SS10[19][10] = 4'h0;
    SS10[20][10] = 4'h0;
    SS10[21][10] = 4'h0;
    SS10[22][10] = 4'h0;
    SS10[23][10] = 4'h0;
    SS10[24][10] = 4'hD;
    SS10[25][10] = 4'hD;
    SS10[26][10] = 4'hD;
    SS10[27][10] = 4'hE;
    SS10[28][10] = 4'hE;
    SS10[29][10] = 4'hE;
    SS10[30][10] = 4'hE;
    SS10[31][10] = 4'hE;
    SS10[32][10] = 4'hE;
    SS10[33][10] = 4'h0;
    SS10[34][10] = 4'h0;
    SS10[35][10] = 4'h0;
    SS10[36][10] = 4'h0;
    SS10[37][10] = 4'h0;
    SS10[38][10] = 4'h0;
    SS10[39][10] = 4'hC;
    SS10[40][10] = 4'hC;
    SS10[41][10] = 4'hC;
    SS10[42][10] = 4'hC;
    SS10[43][10] = 4'hC;
    SS10[44][10] = 4'hC;
    SS10[45][10] = 4'hD;
    SS10[46][10] = 4'hD;
    SS10[47][10] = 4'hD;
    SS10[0][11] = 4'h0;
    SS10[1][11] = 4'h0;
    SS10[2][11] = 4'h0;
    SS10[3][11] = 4'h0;
    SS10[4][11] = 4'h0;
    SS10[5][11] = 4'h0;
    SS10[6][11] = 4'h0;
    SS10[7][11] = 4'h0;
    SS10[8][11] = 4'h0;
    SS10[9][11] = 4'h0;
    SS10[10][11] = 4'h0;
    SS10[11][11] = 4'h0;
    SS10[12][11] = 4'h0;
    SS10[13][11] = 4'h0;
    SS10[14][11] = 4'h0;
    SS10[15][11] = 4'h0;
    SS10[16][11] = 4'h0;
    SS10[17][11] = 4'h0;
    SS10[18][11] = 4'h0;
    SS10[19][11] = 4'h0;
    SS10[20][11] = 4'h0;
    SS10[21][11] = 4'h0;
    SS10[22][11] = 4'h0;
    SS10[23][11] = 4'h0;
    SS10[24][11] = 4'hD;
    SS10[25][11] = 4'hD;
    SS10[26][11] = 4'hD;
    SS10[27][11] = 4'hE;
    SS10[28][11] = 4'hE;
    SS10[29][11] = 4'hE;
    SS10[30][11] = 4'hE;
    SS10[31][11] = 4'hE;
    SS10[32][11] = 4'hE;
    SS10[33][11] = 4'h0;
    SS10[34][11] = 4'h0;
    SS10[35][11] = 4'h0;
    SS10[36][11] = 4'h0;
    SS10[37][11] = 4'h0;
    SS10[38][11] = 4'h0;
    SS10[39][11] = 4'hC;
    SS10[40][11] = 4'hC;
    SS10[41][11] = 4'hC;
    SS10[42][11] = 4'hC;
    SS10[43][11] = 4'hC;
    SS10[44][11] = 4'hC;
    SS10[45][11] = 4'hD;
    SS10[46][11] = 4'hD;
    SS10[47][11] = 4'hD;
    SS10[0][12] = 4'h0;
    SS10[1][12] = 4'h0;
    SS10[2][12] = 4'h0;
    SS10[3][12] = 4'h0;
    SS10[4][12] = 4'h0;
    SS10[5][12] = 4'h0;
    SS10[6][12] = 4'h0;
    SS10[7][12] = 4'h0;
    SS10[8][12] = 4'h0;
    SS10[9][12] = 4'h0;
    SS10[10][12] = 4'h0;
    SS10[11][12] = 4'h0;
    SS10[12][12] = 4'h0;
    SS10[13][12] = 4'h0;
    SS10[14][12] = 4'h0;
    SS10[15][12] = 4'h0;
    SS10[16][12] = 4'h0;
    SS10[17][12] = 4'h0;
    SS10[18][12] = 4'h3;
    SS10[19][12] = 4'h3;
    SS10[20][12] = 4'h3;
    SS10[21][12] = 4'hD;
    SS10[22][12] = 4'hD;
    SS10[23][12] = 4'hD;
    SS10[24][12] = 4'hD;
    SS10[25][12] = 4'hD;
    SS10[26][12] = 4'hD;
    SS10[27][12] = 4'hE;
    SS10[28][12] = 4'hE;
    SS10[29][12] = 4'hE;
    SS10[30][12] = 4'hC;
    SS10[31][12] = 4'hC;
    SS10[32][12] = 4'hC;
    SS10[33][12] = 4'hC;
    SS10[34][12] = 4'hC;
    SS10[35][12] = 4'hC;
    SS10[36][12] = 4'hC;
    SS10[37][12] = 4'hC;
    SS10[38][12] = 4'hC;
    SS10[39][12] = 4'hC;
    SS10[40][12] = 4'hC;
    SS10[41][12] = 4'hC;
    SS10[42][12] = 4'hD;
    SS10[43][12] = 4'hD;
    SS10[44][12] = 4'hD;
    SS10[45][12] = 4'h0;
    SS10[46][12] = 4'h0;
    SS10[47][12] = 4'h0;
    SS10[0][13] = 4'h0;
    SS10[1][13] = 4'h0;
    SS10[2][13] = 4'h0;
    SS10[3][13] = 4'h0;
    SS10[4][13] = 4'h0;
    SS10[5][13] = 4'h0;
    SS10[6][13] = 4'h0;
    SS10[7][13] = 4'h0;
    SS10[8][13] = 4'h0;
    SS10[9][13] = 4'h0;
    SS10[10][13] = 4'h0;
    SS10[11][13] = 4'h0;
    SS10[12][13] = 4'h0;
    SS10[13][13] = 4'h0;
    SS10[14][13] = 4'h0;
    SS10[15][13] = 4'h0;
    SS10[16][13] = 4'h0;
    SS10[17][13] = 4'h0;
    SS10[18][13] = 4'h3;
    SS10[19][13] = 4'h3;
    SS10[20][13] = 4'h3;
    SS10[21][13] = 4'hD;
    SS10[22][13] = 4'hD;
    SS10[23][13] = 4'hD;
    SS10[24][13] = 4'hD;
    SS10[25][13] = 4'hD;
    SS10[26][13] = 4'hD;
    SS10[27][13] = 4'hE;
    SS10[28][13] = 4'hE;
    SS10[29][13] = 4'hE;
    SS10[30][13] = 4'hC;
    SS10[31][13] = 4'hC;
    SS10[32][13] = 4'hC;
    SS10[33][13] = 4'hC;
    SS10[34][13] = 4'hC;
    SS10[35][13] = 4'hC;
    SS10[36][13] = 4'hC;
    SS10[37][13] = 4'hC;
    SS10[38][13] = 4'hC;
    SS10[39][13] = 4'hC;
    SS10[40][13] = 4'hC;
    SS10[41][13] = 4'hC;
    SS10[42][13] = 4'hD;
    SS10[43][13] = 4'hD;
    SS10[44][13] = 4'hD;
    SS10[45][13] = 4'h0;
    SS10[46][13] = 4'h0;
    SS10[47][13] = 4'h0;
    SS10[0][14] = 4'h0;
    SS10[1][14] = 4'h0;
    SS10[2][14] = 4'h0;
    SS10[3][14] = 4'h0;
    SS10[4][14] = 4'h0;
    SS10[5][14] = 4'h0;
    SS10[6][14] = 4'h0;
    SS10[7][14] = 4'h0;
    SS10[8][14] = 4'h0;
    SS10[9][14] = 4'h0;
    SS10[10][14] = 4'h0;
    SS10[11][14] = 4'h0;
    SS10[12][14] = 4'h0;
    SS10[13][14] = 4'h0;
    SS10[14][14] = 4'h0;
    SS10[15][14] = 4'h0;
    SS10[16][14] = 4'h0;
    SS10[17][14] = 4'h0;
    SS10[18][14] = 4'h3;
    SS10[19][14] = 4'h3;
    SS10[20][14] = 4'h3;
    SS10[21][14] = 4'hD;
    SS10[22][14] = 4'hD;
    SS10[23][14] = 4'hD;
    SS10[24][14] = 4'hD;
    SS10[25][14] = 4'hD;
    SS10[26][14] = 4'hD;
    SS10[27][14] = 4'hE;
    SS10[28][14] = 4'hE;
    SS10[29][14] = 4'hE;
    SS10[30][14] = 4'hC;
    SS10[31][14] = 4'hC;
    SS10[32][14] = 4'hC;
    SS10[33][14] = 4'hC;
    SS10[34][14] = 4'hC;
    SS10[35][14] = 4'hC;
    SS10[36][14] = 4'hC;
    SS10[37][14] = 4'hC;
    SS10[38][14] = 4'hC;
    SS10[39][14] = 4'hC;
    SS10[40][14] = 4'hC;
    SS10[41][14] = 4'hC;
    SS10[42][14] = 4'hD;
    SS10[43][14] = 4'hD;
    SS10[44][14] = 4'hD;
    SS10[45][14] = 4'h0;
    SS10[46][14] = 4'h0;
    SS10[47][14] = 4'h0;
    SS10[0][15] = 4'h0;
    SS10[1][15] = 4'h0;
    SS10[2][15] = 4'h0;
    SS10[3][15] = 4'h0;
    SS10[4][15] = 4'h0;
    SS10[5][15] = 4'h0;
    SS10[6][15] = 4'h0;
    SS10[7][15] = 4'h0;
    SS10[8][15] = 4'h0;
    SS10[9][15] = 4'h0;
    SS10[10][15] = 4'h0;
    SS10[11][15] = 4'h0;
    SS10[12][15] = 4'h0;
    SS10[13][15] = 4'h0;
    SS10[14][15] = 4'h0;
    SS10[15][15] = 4'h0;
    SS10[16][15] = 4'h0;
    SS10[17][15] = 4'h0;
    SS10[18][15] = 4'hD;
    SS10[19][15] = 4'hD;
    SS10[20][15] = 4'hD;
    SS10[21][15] = 4'hD;
    SS10[22][15] = 4'hD;
    SS10[23][15] = 4'hD;
    SS10[24][15] = 4'hE;
    SS10[25][15] = 4'hE;
    SS10[26][15] = 4'hE;
    SS10[27][15] = 4'hC;
    SS10[28][15] = 4'hC;
    SS10[29][15] = 4'hC;
    SS10[30][15] = 4'hC;
    SS10[31][15] = 4'hC;
    SS10[32][15] = 4'hC;
    SS10[33][15] = 4'hC;
    SS10[34][15] = 4'hC;
    SS10[35][15] = 4'hC;
    SS10[36][15] = 4'hD;
    SS10[37][15] = 4'hD;
    SS10[38][15] = 4'hD;
    SS10[39][15] = 4'hE;
    SS10[40][15] = 4'hE;
    SS10[41][15] = 4'hE;
    SS10[42][15] = 4'h0;
    SS10[43][15] = 4'h0;
    SS10[44][15] = 4'h0;
    SS10[45][15] = 4'h0;
    SS10[46][15] = 4'h0;
    SS10[47][15] = 4'h0;
    SS10[0][16] = 4'h0;
    SS10[1][16] = 4'h0;
    SS10[2][16] = 4'h0;
    SS10[3][16] = 4'h0;
    SS10[4][16] = 4'h0;
    SS10[5][16] = 4'h0;
    SS10[6][16] = 4'h0;
    SS10[7][16] = 4'h0;
    SS10[8][16] = 4'h0;
    SS10[9][16] = 4'h0;
    SS10[10][16] = 4'h0;
    SS10[11][16] = 4'h0;
    SS10[12][16] = 4'h0;
    SS10[13][16] = 4'h0;
    SS10[14][16] = 4'h0;
    SS10[15][16] = 4'h0;
    SS10[16][16] = 4'h0;
    SS10[17][16] = 4'h0;
    SS10[18][16] = 4'hD;
    SS10[19][16] = 4'hD;
    SS10[20][16] = 4'hD;
    SS10[21][16] = 4'hD;
    SS10[22][16] = 4'hD;
    SS10[23][16] = 4'hD;
    SS10[24][16] = 4'hE;
    SS10[25][16] = 4'hE;
    SS10[26][16] = 4'hE;
    SS10[27][16] = 4'hC;
    SS10[28][16] = 4'hC;
    SS10[29][16] = 4'hC;
    SS10[30][16] = 4'hC;
    SS10[31][16] = 4'hC;
    SS10[32][16] = 4'hC;
    SS10[33][16] = 4'hC;
    SS10[34][16] = 4'hC;
    SS10[35][16] = 4'hC;
    SS10[36][16] = 4'hD;
    SS10[37][16] = 4'hD;
    SS10[38][16] = 4'hD;
    SS10[39][16] = 4'hE;
    SS10[40][16] = 4'hE;
    SS10[41][16] = 4'hE;
    SS10[42][16] = 4'h0;
    SS10[43][16] = 4'h0;
    SS10[44][16] = 4'h0;
    SS10[45][16] = 4'h0;
    SS10[46][16] = 4'h0;
    SS10[47][16] = 4'h0;
    SS10[0][17] = 4'h0;
    SS10[1][17] = 4'h0;
    SS10[2][17] = 4'h0;
    SS10[3][17] = 4'h0;
    SS10[4][17] = 4'h0;
    SS10[5][17] = 4'h0;
    SS10[6][17] = 4'h0;
    SS10[7][17] = 4'h0;
    SS10[8][17] = 4'h0;
    SS10[9][17] = 4'h0;
    SS10[10][17] = 4'h0;
    SS10[11][17] = 4'h0;
    SS10[12][17] = 4'h0;
    SS10[13][17] = 4'h0;
    SS10[14][17] = 4'h0;
    SS10[15][17] = 4'h0;
    SS10[16][17] = 4'h0;
    SS10[17][17] = 4'h0;
    SS10[18][17] = 4'hD;
    SS10[19][17] = 4'hD;
    SS10[20][17] = 4'hD;
    SS10[21][17] = 4'hD;
    SS10[22][17] = 4'hD;
    SS10[23][17] = 4'hD;
    SS10[24][17] = 4'hE;
    SS10[25][17] = 4'hE;
    SS10[26][17] = 4'hE;
    SS10[27][17] = 4'hC;
    SS10[28][17] = 4'hC;
    SS10[29][17] = 4'hC;
    SS10[30][17] = 4'hC;
    SS10[31][17] = 4'hC;
    SS10[32][17] = 4'hC;
    SS10[33][17] = 4'hC;
    SS10[34][17] = 4'hC;
    SS10[35][17] = 4'hC;
    SS10[36][17] = 4'hD;
    SS10[37][17] = 4'hD;
    SS10[38][17] = 4'hD;
    SS10[39][17] = 4'hE;
    SS10[40][17] = 4'hE;
    SS10[41][17] = 4'hE;
    SS10[42][17] = 4'h0;
    SS10[43][17] = 4'h0;
    SS10[44][17] = 4'h0;
    SS10[45][17] = 4'h0;
    SS10[46][17] = 4'h0;
    SS10[47][17] = 4'h0;
    SS10[0][18] = 4'h0;
    SS10[1][18] = 4'h0;
    SS10[2][18] = 4'h0;
    SS10[3][18] = 4'h0;
    SS10[4][18] = 4'h0;
    SS10[5][18] = 4'h0;
    SS10[6][18] = 4'hD;
    SS10[7][18] = 4'hD;
    SS10[8][18] = 4'hD;
    SS10[9][18] = 4'hD;
    SS10[10][18] = 4'hD;
    SS10[11][18] = 4'hD;
    SS10[12][18] = 4'hD;
    SS10[13][18] = 4'hD;
    SS10[14][18] = 4'hD;
    SS10[15][18] = 4'hC;
    SS10[16][18] = 4'hC;
    SS10[17][18] = 4'hC;
    SS10[18][18] = 4'hD;
    SS10[19][18] = 4'hD;
    SS10[20][18] = 4'hD;
    SS10[21][18] = 4'hC;
    SS10[22][18] = 4'hC;
    SS10[23][18] = 4'hC;
    SS10[24][18] = 4'hC;
    SS10[25][18] = 4'hC;
    SS10[26][18] = 4'hC;
    SS10[27][18] = 4'hC;
    SS10[28][18] = 4'hC;
    SS10[29][18] = 4'hC;
    SS10[30][18] = 4'hC;
    SS10[31][18] = 4'hC;
    SS10[32][18] = 4'hC;
    SS10[33][18] = 4'hD;
    SS10[34][18] = 4'hD;
    SS10[35][18] = 4'hD;
    SS10[36][18] = 4'hE;
    SS10[37][18] = 4'hE;
    SS10[38][18] = 4'hE;
    SS10[39][18] = 4'h0;
    SS10[40][18] = 4'h0;
    SS10[41][18] = 4'h0;
    SS10[42][18] = 4'h0;
    SS10[43][18] = 4'h0;
    SS10[44][18] = 4'h0;
    SS10[45][18] = 4'h0;
    SS10[46][18] = 4'h0;
    SS10[47][18] = 4'h0;
    SS10[0][19] = 4'h0;
    SS10[1][19] = 4'h0;
    SS10[2][19] = 4'h0;
    SS10[3][19] = 4'h0;
    SS10[4][19] = 4'h0;
    SS10[5][19] = 4'h0;
    SS10[6][19] = 4'hD;
    SS10[7][19] = 4'hD;
    SS10[8][19] = 4'hD;
    SS10[9][19] = 4'hD;
    SS10[10][19] = 4'hD;
    SS10[11][19] = 4'hD;
    SS10[12][19] = 4'hD;
    SS10[13][19] = 4'hD;
    SS10[14][19] = 4'hD;
    SS10[15][19] = 4'hC;
    SS10[16][19] = 4'hC;
    SS10[17][19] = 4'hC;
    SS10[18][19] = 4'hD;
    SS10[19][19] = 4'hD;
    SS10[20][19] = 4'hD;
    SS10[21][19] = 4'hC;
    SS10[22][19] = 4'hC;
    SS10[23][19] = 4'hC;
    SS10[24][19] = 4'hC;
    SS10[25][19] = 4'hC;
    SS10[26][19] = 4'hC;
    SS10[27][19] = 4'hC;
    SS10[28][19] = 4'hC;
    SS10[29][19] = 4'hC;
    SS10[30][19] = 4'hC;
    SS10[31][19] = 4'hC;
    SS10[32][19] = 4'hC;
    SS10[33][19] = 4'hD;
    SS10[34][19] = 4'hD;
    SS10[35][19] = 4'hD;
    SS10[36][19] = 4'hE;
    SS10[37][19] = 4'hE;
    SS10[38][19] = 4'hE;
    SS10[39][19] = 4'h0;
    SS10[40][19] = 4'h0;
    SS10[41][19] = 4'h0;
    SS10[42][19] = 4'h0;
    SS10[43][19] = 4'h0;
    SS10[44][19] = 4'h0;
    SS10[45][19] = 4'h0;
    SS10[46][19] = 4'h0;
    SS10[47][19] = 4'h0;
    SS10[0][20] = 4'h0;
    SS10[1][20] = 4'h0;
    SS10[2][20] = 4'h0;
    SS10[3][20] = 4'h0;
    SS10[4][20] = 4'h0;
    SS10[5][20] = 4'h0;
    SS10[6][20] = 4'hD;
    SS10[7][20] = 4'hD;
    SS10[8][20] = 4'hD;
    SS10[9][20] = 4'hD;
    SS10[10][20] = 4'hD;
    SS10[11][20] = 4'hD;
    SS10[12][20] = 4'hD;
    SS10[13][20] = 4'hD;
    SS10[14][20] = 4'hD;
    SS10[15][20] = 4'hC;
    SS10[16][20] = 4'hC;
    SS10[17][20] = 4'hC;
    SS10[18][20] = 4'hD;
    SS10[19][20] = 4'hD;
    SS10[20][20] = 4'hD;
    SS10[21][20] = 4'hC;
    SS10[22][20] = 4'hC;
    SS10[23][20] = 4'hC;
    SS10[24][20] = 4'hC;
    SS10[25][20] = 4'hC;
    SS10[26][20] = 4'hC;
    SS10[27][20] = 4'hC;
    SS10[28][20] = 4'hC;
    SS10[29][20] = 4'hC;
    SS10[30][20] = 4'hC;
    SS10[31][20] = 4'hC;
    SS10[32][20] = 4'hC;
    SS10[33][20] = 4'hD;
    SS10[34][20] = 4'hD;
    SS10[35][20] = 4'hD;
    SS10[36][20] = 4'hE;
    SS10[37][20] = 4'hE;
    SS10[38][20] = 4'hE;
    SS10[39][20] = 4'h0;
    SS10[40][20] = 4'h0;
    SS10[41][20] = 4'h0;
    SS10[42][20] = 4'h0;
    SS10[43][20] = 4'h0;
    SS10[44][20] = 4'h0;
    SS10[45][20] = 4'h0;
    SS10[46][20] = 4'h0;
    SS10[47][20] = 4'h0;
    SS10[0][21] = 4'hC;
    SS10[1][21] = 4'hC;
    SS10[2][21] = 4'hC;
    SS10[3][21] = 4'hC;
    SS10[4][21] = 4'hC;
    SS10[5][21] = 4'hC;
    SS10[6][21] = 4'hC;
    SS10[7][21] = 4'hC;
    SS10[8][21] = 4'hC;
    SS10[9][21] = 4'hC;
    SS10[10][21] = 4'hC;
    SS10[11][21] = 4'hC;
    SS10[12][21] = 4'hC;
    SS10[13][21] = 4'hC;
    SS10[14][21] = 4'hC;
    SS10[15][21] = 4'hC;
    SS10[16][21] = 4'hC;
    SS10[17][21] = 4'hC;
    SS10[18][21] = 4'hA;
    SS10[19][21] = 4'hA;
    SS10[20][21] = 4'hA;
    SS10[21][21] = 4'hD;
    SS10[22][21] = 4'hD;
    SS10[23][21] = 4'hD;
    SS10[24][21] = 4'hC;
    SS10[25][21] = 4'hC;
    SS10[26][21] = 4'hC;
    SS10[27][21] = 4'hD;
    SS10[28][21] = 4'hD;
    SS10[29][21] = 4'hD;
    SS10[30][21] = 4'hE;
    SS10[31][21] = 4'hE;
    SS10[32][21] = 4'hE;
    SS10[33][21] = 4'hE;
    SS10[34][21] = 4'hE;
    SS10[35][21] = 4'hE;
    SS10[36][21] = 4'h0;
    SS10[37][21] = 4'h0;
    SS10[38][21] = 4'h0;
    SS10[39][21] = 4'h0;
    SS10[40][21] = 4'h0;
    SS10[41][21] = 4'h0;
    SS10[42][21] = 4'h0;
    SS10[43][21] = 4'h0;
    SS10[44][21] = 4'h0;
    SS10[45][21] = 4'h0;
    SS10[46][21] = 4'h0;
    SS10[47][21] = 4'h0;
    SS10[0][22] = 4'hC;
    SS10[1][22] = 4'hC;
    SS10[2][22] = 4'hC;
    SS10[3][22] = 4'hC;
    SS10[4][22] = 4'hC;
    SS10[5][22] = 4'hC;
    SS10[6][22] = 4'hC;
    SS10[7][22] = 4'hC;
    SS10[8][22] = 4'hC;
    SS10[9][22] = 4'hC;
    SS10[10][22] = 4'hC;
    SS10[11][22] = 4'hC;
    SS10[12][22] = 4'hC;
    SS10[13][22] = 4'hC;
    SS10[14][22] = 4'hC;
    SS10[15][22] = 4'hC;
    SS10[16][22] = 4'hC;
    SS10[17][22] = 4'hC;
    SS10[18][22] = 4'hA;
    SS10[19][22] = 4'hA;
    SS10[20][22] = 4'hA;
    SS10[21][22] = 4'hD;
    SS10[22][22] = 4'hD;
    SS10[23][22] = 4'hD;
    SS10[24][22] = 4'hC;
    SS10[25][22] = 4'hC;
    SS10[26][22] = 4'hC;
    SS10[27][22] = 4'hD;
    SS10[28][22] = 4'hD;
    SS10[29][22] = 4'hD;
    SS10[30][22] = 4'hE;
    SS10[31][22] = 4'hE;
    SS10[32][22] = 4'hE;
    SS10[33][22] = 4'hE;
    SS10[34][22] = 4'hE;
    SS10[35][22] = 4'hE;
    SS10[36][22] = 4'h0;
    SS10[37][22] = 4'h0;
    SS10[38][22] = 4'h0;
    SS10[39][22] = 4'h0;
    SS10[40][22] = 4'h0;
    SS10[41][22] = 4'h0;
    SS10[42][22] = 4'h0;
    SS10[43][22] = 4'h0;
    SS10[44][22] = 4'h0;
    SS10[45][22] = 4'h0;
    SS10[46][22] = 4'h0;
    SS10[47][22] = 4'h0;
    SS10[0][23] = 4'hC;
    SS10[1][23] = 4'hC;
    SS10[2][23] = 4'hC;
    SS10[3][23] = 4'hC;
    SS10[4][23] = 4'hC;
    SS10[5][23] = 4'hC;
    SS10[6][23] = 4'hC;
    SS10[7][23] = 4'hC;
    SS10[8][23] = 4'hC;
    SS10[9][23] = 4'hC;
    SS10[10][23] = 4'hC;
    SS10[11][23] = 4'hC;
    SS10[12][23] = 4'hC;
    SS10[13][23] = 4'hC;
    SS10[14][23] = 4'hC;
    SS10[15][23] = 4'hC;
    SS10[16][23] = 4'hC;
    SS10[17][23] = 4'hC;
    SS10[18][23] = 4'hA;
    SS10[19][23] = 4'hA;
    SS10[20][23] = 4'hA;
    SS10[21][23] = 4'hD;
    SS10[22][23] = 4'hD;
    SS10[23][23] = 4'hD;
    SS10[24][23] = 4'hC;
    SS10[25][23] = 4'hC;
    SS10[26][23] = 4'hC;
    SS10[27][23] = 4'hD;
    SS10[28][23] = 4'hD;
    SS10[29][23] = 4'hD;
    SS10[30][23] = 4'hE;
    SS10[31][23] = 4'hE;
    SS10[32][23] = 4'hE;
    SS10[33][23] = 4'hE;
    SS10[34][23] = 4'hE;
    SS10[35][23] = 4'hE;
    SS10[36][23] = 4'h0;
    SS10[37][23] = 4'h0;
    SS10[38][23] = 4'h0;
    SS10[39][23] = 4'h0;
    SS10[40][23] = 4'h0;
    SS10[41][23] = 4'h0;
    SS10[42][23] = 4'h0;
    SS10[43][23] = 4'h0;
    SS10[44][23] = 4'h0;
    SS10[45][23] = 4'h0;
    SS10[46][23] = 4'h0;
    SS10[47][23] = 4'h0;
    SS10[0][24] = 4'hC;
    SS10[1][24] = 4'hC;
    SS10[2][24] = 4'hC;
    SS10[3][24] = 4'hC;
    SS10[4][24] = 4'hC;
    SS10[5][24] = 4'hC;
    SS10[6][24] = 4'hC;
    SS10[7][24] = 4'hC;
    SS10[8][24] = 4'hC;
    SS10[9][24] = 4'hC;
    SS10[10][24] = 4'hC;
    SS10[11][24] = 4'hC;
    SS10[12][24] = 4'hC;
    SS10[13][24] = 4'hC;
    SS10[14][24] = 4'hC;
    SS10[15][24] = 4'hC;
    SS10[16][24] = 4'hC;
    SS10[17][24] = 4'hC;
    SS10[18][24] = 4'hA;
    SS10[19][24] = 4'hA;
    SS10[20][24] = 4'hA;
    SS10[21][24] = 4'hD;
    SS10[22][24] = 4'hD;
    SS10[23][24] = 4'hD;
    SS10[24][24] = 4'hC;
    SS10[25][24] = 4'hC;
    SS10[26][24] = 4'hC;
    SS10[27][24] = 4'hD;
    SS10[28][24] = 4'hD;
    SS10[29][24] = 4'hD;
    SS10[30][24] = 4'hE;
    SS10[31][24] = 4'hE;
    SS10[32][24] = 4'hE;
    SS10[33][24] = 4'hE;
    SS10[34][24] = 4'hE;
    SS10[35][24] = 4'hE;
    SS10[36][24] = 4'h0;
    SS10[37][24] = 4'h0;
    SS10[38][24] = 4'h0;
    SS10[39][24] = 4'h0;
    SS10[40][24] = 4'h0;
    SS10[41][24] = 4'h0;
    SS10[42][24] = 4'h0;
    SS10[43][24] = 4'h0;
    SS10[44][24] = 4'h0;
    SS10[45][24] = 4'h0;
    SS10[46][24] = 4'h0;
    SS10[47][24] = 4'h0;
    SS10[0][25] = 4'hC;
    SS10[1][25] = 4'hC;
    SS10[2][25] = 4'hC;
    SS10[3][25] = 4'hC;
    SS10[4][25] = 4'hC;
    SS10[5][25] = 4'hC;
    SS10[6][25] = 4'hC;
    SS10[7][25] = 4'hC;
    SS10[8][25] = 4'hC;
    SS10[9][25] = 4'hC;
    SS10[10][25] = 4'hC;
    SS10[11][25] = 4'hC;
    SS10[12][25] = 4'hC;
    SS10[13][25] = 4'hC;
    SS10[14][25] = 4'hC;
    SS10[15][25] = 4'hC;
    SS10[16][25] = 4'hC;
    SS10[17][25] = 4'hC;
    SS10[18][25] = 4'hA;
    SS10[19][25] = 4'hA;
    SS10[20][25] = 4'hA;
    SS10[21][25] = 4'hD;
    SS10[22][25] = 4'hD;
    SS10[23][25] = 4'hD;
    SS10[24][25] = 4'hC;
    SS10[25][25] = 4'hC;
    SS10[26][25] = 4'hC;
    SS10[27][25] = 4'hD;
    SS10[28][25] = 4'hD;
    SS10[29][25] = 4'hD;
    SS10[30][25] = 4'hE;
    SS10[31][25] = 4'hE;
    SS10[32][25] = 4'hE;
    SS10[33][25] = 4'hE;
    SS10[34][25] = 4'hE;
    SS10[35][25] = 4'hE;
    SS10[36][25] = 4'h0;
    SS10[37][25] = 4'h0;
    SS10[38][25] = 4'h0;
    SS10[39][25] = 4'h0;
    SS10[40][25] = 4'h0;
    SS10[41][25] = 4'h0;
    SS10[42][25] = 4'h0;
    SS10[43][25] = 4'h0;
    SS10[44][25] = 4'h0;
    SS10[45][25] = 4'h0;
    SS10[46][25] = 4'h0;
    SS10[47][25] = 4'h0;
    SS10[0][26] = 4'hC;
    SS10[1][26] = 4'hC;
    SS10[2][26] = 4'hC;
    SS10[3][26] = 4'hC;
    SS10[4][26] = 4'hC;
    SS10[5][26] = 4'hC;
    SS10[6][26] = 4'hC;
    SS10[7][26] = 4'hC;
    SS10[8][26] = 4'hC;
    SS10[9][26] = 4'hC;
    SS10[10][26] = 4'hC;
    SS10[11][26] = 4'hC;
    SS10[12][26] = 4'hC;
    SS10[13][26] = 4'hC;
    SS10[14][26] = 4'hC;
    SS10[15][26] = 4'hC;
    SS10[16][26] = 4'hC;
    SS10[17][26] = 4'hC;
    SS10[18][26] = 4'hA;
    SS10[19][26] = 4'hA;
    SS10[20][26] = 4'hA;
    SS10[21][26] = 4'hD;
    SS10[22][26] = 4'hD;
    SS10[23][26] = 4'hD;
    SS10[24][26] = 4'hC;
    SS10[25][26] = 4'hC;
    SS10[26][26] = 4'hC;
    SS10[27][26] = 4'hD;
    SS10[28][26] = 4'hD;
    SS10[29][26] = 4'hD;
    SS10[30][26] = 4'hE;
    SS10[31][26] = 4'hE;
    SS10[32][26] = 4'hE;
    SS10[33][26] = 4'hE;
    SS10[34][26] = 4'hE;
    SS10[35][26] = 4'hE;
    SS10[36][26] = 4'h0;
    SS10[37][26] = 4'h0;
    SS10[38][26] = 4'h0;
    SS10[39][26] = 4'h0;
    SS10[40][26] = 4'h0;
    SS10[41][26] = 4'h0;
    SS10[42][26] = 4'h0;
    SS10[43][26] = 4'h0;
    SS10[44][26] = 4'h0;
    SS10[45][26] = 4'h0;
    SS10[46][26] = 4'h0;
    SS10[47][26] = 4'h0;
    SS10[0][27] = 4'h0;
    SS10[1][27] = 4'h0;
    SS10[2][27] = 4'h0;
    SS10[3][27] = 4'h0;
    SS10[4][27] = 4'h0;
    SS10[5][27] = 4'h0;
    SS10[6][27] = 4'hD;
    SS10[7][27] = 4'hD;
    SS10[8][27] = 4'hD;
    SS10[9][27] = 4'hD;
    SS10[10][27] = 4'hD;
    SS10[11][27] = 4'hD;
    SS10[12][27] = 4'hD;
    SS10[13][27] = 4'hD;
    SS10[14][27] = 4'hD;
    SS10[15][27] = 4'hC;
    SS10[16][27] = 4'hC;
    SS10[17][27] = 4'hC;
    SS10[18][27] = 4'hD;
    SS10[19][27] = 4'hD;
    SS10[20][27] = 4'hD;
    SS10[21][27] = 4'hC;
    SS10[22][27] = 4'hC;
    SS10[23][27] = 4'hC;
    SS10[24][27] = 4'hC;
    SS10[25][27] = 4'hC;
    SS10[26][27] = 4'hC;
    SS10[27][27] = 4'hC;
    SS10[28][27] = 4'hC;
    SS10[29][27] = 4'hC;
    SS10[30][27] = 4'hC;
    SS10[31][27] = 4'hC;
    SS10[32][27] = 4'hC;
    SS10[33][27] = 4'hD;
    SS10[34][27] = 4'hD;
    SS10[35][27] = 4'hD;
    SS10[36][27] = 4'hE;
    SS10[37][27] = 4'hE;
    SS10[38][27] = 4'hE;
    SS10[39][27] = 4'h0;
    SS10[40][27] = 4'h0;
    SS10[41][27] = 4'h0;
    SS10[42][27] = 4'h0;
    SS10[43][27] = 4'h0;
    SS10[44][27] = 4'h0;
    SS10[45][27] = 4'h0;
    SS10[46][27] = 4'h0;
    SS10[47][27] = 4'h0;
    SS10[0][28] = 4'h0;
    SS10[1][28] = 4'h0;
    SS10[2][28] = 4'h0;
    SS10[3][28] = 4'h0;
    SS10[4][28] = 4'h0;
    SS10[5][28] = 4'h0;
    SS10[6][28] = 4'hD;
    SS10[7][28] = 4'hD;
    SS10[8][28] = 4'hD;
    SS10[9][28] = 4'hD;
    SS10[10][28] = 4'hD;
    SS10[11][28] = 4'hD;
    SS10[12][28] = 4'hD;
    SS10[13][28] = 4'hD;
    SS10[14][28] = 4'hD;
    SS10[15][28] = 4'hC;
    SS10[16][28] = 4'hC;
    SS10[17][28] = 4'hC;
    SS10[18][28] = 4'hD;
    SS10[19][28] = 4'hD;
    SS10[20][28] = 4'hD;
    SS10[21][28] = 4'hC;
    SS10[22][28] = 4'hC;
    SS10[23][28] = 4'hC;
    SS10[24][28] = 4'hC;
    SS10[25][28] = 4'hC;
    SS10[26][28] = 4'hC;
    SS10[27][28] = 4'hC;
    SS10[28][28] = 4'hC;
    SS10[29][28] = 4'hC;
    SS10[30][28] = 4'hC;
    SS10[31][28] = 4'hC;
    SS10[32][28] = 4'hC;
    SS10[33][28] = 4'hD;
    SS10[34][28] = 4'hD;
    SS10[35][28] = 4'hD;
    SS10[36][28] = 4'hE;
    SS10[37][28] = 4'hE;
    SS10[38][28] = 4'hE;
    SS10[39][28] = 4'h0;
    SS10[40][28] = 4'h0;
    SS10[41][28] = 4'h0;
    SS10[42][28] = 4'h0;
    SS10[43][28] = 4'h0;
    SS10[44][28] = 4'h0;
    SS10[45][28] = 4'h0;
    SS10[46][28] = 4'h0;
    SS10[47][28] = 4'h0;
    SS10[0][29] = 4'h0;
    SS10[1][29] = 4'h0;
    SS10[2][29] = 4'h0;
    SS10[3][29] = 4'h0;
    SS10[4][29] = 4'h0;
    SS10[5][29] = 4'h0;
    SS10[6][29] = 4'hD;
    SS10[7][29] = 4'hD;
    SS10[8][29] = 4'hD;
    SS10[9][29] = 4'hD;
    SS10[10][29] = 4'hD;
    SS10[11][29] = 4'hD;
    SS10[12][29] = 4'hD;
    SS10[13][29] = 4'hD;
    SS10[14][29] = 4'hD;
    SS10[15][29] = 4'hC;
    SS10[16][29] = 4'hC;
    SS10[17][29] = 4'hC;
    SS10[18][29] = 4'hD;
    SS10[19][29] = 4'hD;
    SS10[20][29] = 4'hD;
    SS10[21][29] = 4'hC;
    SS10[22][29] = 4'hC;
    SS10[23][29] = 4'hC;
    SS10[24][29] = 4'hC;
    SS10[25][29] = 4'hC;
    SS10[26][29] = 4'hC;
    SS10[27][29] = 4'hC;
    SS10[28][29] = 4'hC;
    SS10[29][29] = 4'hC;
    SS10[30][29] = 4'hC;
    SS10[31][29] = 4'hC;
    SS10[32][29] = 4'hC;
    SS10[33][29] = 4'hD;
    SS10[34][29] = 4'hD;
    SS10[35][29] = 4'hD;
    SS10[36][29] = 4'hE;
    SS10[37][29] = 4'hE;
    SS10[38][29] = 4'hE;
    SS10[39][29] = 4'h0;
    SS10[40][29] = 4'h0;
    SS10[41][29] = 4'h0;
    SS10[42][29] = 4'h0;
    SS10[43][29] = 4'h0;
    SS10[44][29] = 4'h0;
    SS10[45][29] = 4'h0;
    SS10[46][29] = 4'h0;
    SS10[47][29] = 4'h0;
    SS10[0][30] = 4'h0;
    SS10[1][30] = 4'h0;
    SS10[2][30] = 4'h0;
    SS10[3][30] = 4'h0;
    SS10[4][30] = 4'h0;
    SS10[5][30] = 4'h0;
    SS10[6][30] = 4'h0;
    SS10[7][30] = 4'h0;
    SS10[8][30] = 4'h0;
    SS10[9][30] = 4'h0;
    SS10[10][30] = 4'h0;
    SS10[11][30] = 4'h0;
    SS10[12][30] = 4'h0;
    SS10[13][30] = 4'h0;
    SS10[14][30] = 4'h0;
    SS10[15][30] = 4'h0;
    SS10[16][30] = 4'h0;
    SS10[17][30] = 4'h0;
    SS10[18][30] = 4'hD;
    SS10[19][30] = 4'hD;
    SS10[20][30] = 4'hD;
    SS10[21][30] = 4'hD;
    SS10[22][30] = 4'hD;
    SS10[23][30] = 4'hD;
    SS10[24][30] = 4'hE;
    SS10[25][30] = 4'hE;
    SS10[26][30] = 4'hE;
    SS10[27][30] = 4'hC;
    SS10[28][30] = 4'hC;
    SS10[29][30] = 4'hC;
    SS10[30][30] = 4'hC;
    SS10[31][30] = 4'hC;
    SS10[32][30] = 4'hC;
    SS10[33][30] = 4'hC;
    SS10[34][30] = 4'hC;
    SS10[35][30] = 4'hC;
    SS10[36][30] = 4'hD;
    SS10[37][30] = 4'hD;
    SS10[38][30] = 4'hD;
    SS10[39][30] = 4'hE;
    SS10[40][30] = 4'hE;
    SS10[41][30] = 4'hE;
    SS10[42][30] = 4'h0;
    SS10[43][30] = 4'h0;
    SS10[44][30] = 4'h0;
    SS10[45][30] = 4'h0;
    SS10[46][30] = 4'h0;
    SS10[47][30] = 4'h0;
    SS10[0][31] = 4'h0;
    SS10[1][31] = 4'h0;
    SS10[2][31] = 4'h0;
    SS10[3][31] = 4'h0;
    SS10[4][31] = 4'h0;
    SS10[5][31] = 4'h0;
    SS10[6][31] = 4'h0;
    SS10[7][31] = 4'h0;
    SS10[8][31] = 4'h0;
    SS10[9][31] = 4'h0;
    SS10[10][31] = 4'h0;
    SS10[11][31] = 4'h0;
    SS10[12][31] = 4'h0;
    SS10[13][31] = 4'h0;
    SS10[14][31] = 4'h0;
    SS10[15][31] = 4'h0;
    SS10[16][31] = 4'h0;
    SS10[17][31] = 4'h0;
    SS10[18][31] = 4'hD;
    SS10[19][31] = 4'hD;
    SS10[20][31] = 4'hD;
    SS10[21][31] = 4'hD;
    SS10[22][31] = 4'hD;
    SS10[23][31] = 4'hD;
    SS10[24][31] = 4'hE;
    SS10[25][31] = 4'hE;
    SS10[26][31] = 4'hE;
    SS10[27][31] = 4'hC;
    SS10[28][31] = 4'hC;
    SS10[29][31] = 4'hC;
    SS10[30][31] = 4'hC;
    SS10[31][31] = 4'hC;
    SS10[32][31] = 4'hC;
    SS10[33][31] = 4'hC;
    SS10[34][31] = 4'hC;
    SS10[35][31] = 4'hC;
    SS10[36][31] = 4'hD;
    SS10[37][31] = 4'hD;
    SS10[38][31] = 4'hD;
    SS10[39][31] = 4'hE;
    SS10[40][31] = 4'hE;
    SS10[41][31] = 4'hE;
    SS10[42][31] = 4'h0;
    SS10[43][31] = 4'h0;
    SS10[44][31] = 4'h0;
    SS10[45][31] = 4'h0;
    SS10[46][31] = 4'h0;
    SS10[47][31] = 4'h0;
    SS10[0][32] = 4'h0;
    SS10[1][32] = 4'h0;
    SS10[2][32] = 4'h0;
    SS10[3][32] = 4'h0;
    SS10[4][32] = 4'h0;
    SS10[5][32] = 4'h0;
    SS10[6][32] = 4'h0;
    SS10[7][32] = 4'h0;
    SS10[8][32] = 4'h0;
    SS10[9][32] = 4'h0;
    SS10[10][32] = 4'h0;
    SS10[11][32] = 4'h0;
    SS10[12][32] = 4'h0;
    SS10[13][32] = 4'h0;
    SS10[14][32] = 4'h0;
    SS10[15][32] = 4'h0;
    SS10[16][32] = 4'h0;
    SS10[17][32] = 4'h0;
    SS10[18][32] = 4'hD;
    SS10[19][32] = 4'hD;
    SS10[20][32] = 4'hD;
    SS10[21][32] = 4'hD;
    SS10[22][32] = 4'hD;
    SS10[23][32] = 4'hD;
    SS10[24][32] = 4'hE;
    SS10[25][32] = 4'hE;
    SS10[26][32] = 4'hE;
    SS10[27][32] = 4'hC;
    SS10[28][32] = 4'hC;
    SS10[29][32] = 4'hC;
    SS10[30][32] = 4'hC;
    SS10[31][32] = 4'hC;
    SS10[32][32] = 4'hC;
    SS10[33][32] = 4'hC;
    SS10[34][32] = 4'hC;
    SS10[35][32] = 4'hC;
    SS10[36][32] = 4'hD;
    SS10[37][32] = 4'hD;
    SS10[38][32] = 4'hD;
    SS10[39][32] = 4'hE;
    SS10[40][32] = 4'hE;
    SS10[41][32] = 4'hE;
    SS10[42][32] = 4'h0;
    SS10[43][32] = 4'h0;
    SS10[44][32] = 4'h0;
    SS10[45][32] = 4'h0;
    SS10[46][32] = 4'h0;
    SS10[47][32] = 4'h0;
    SS10[0][33] = 4'h0;
    SS10[1][33] = 4'h0;
    SS10[2][33] = 4'h0;
    SS10[3][33] = 4'h0;
    SS10[4][33] = 4'h0;
    SS10[5][33] = 4'h0;
    SS10[6][33] = 4'h0;
    SS10[7][33] = 4'h0;
    SS10[8][33] = 4'h0;
    SS10[9][33] = 4'h0;
    SS10[10][33] = 4'h0;
    SS10[11][33] = 4'h0;
    SS10[12][33] = 4'h0;
    SS10[13][33] = 4'h0;
    SS10[14][33] = 4'h0;
    SS10[15][33] = 4'h0;
    SS10[16][33] = 4'h0;
    SS10[17][33] = 4'h0;
    SS10[18][33] = 4'h3;
    SS10[19][33] = 4'h3;
    SS10[20][33] = 4'h3;
    SS10[21][33] = 4'hD;
    SS10[22][33] = 4'hD;
    SS10[23][33] = 4'hD;
    SS10[24][33] = 4'hD;
    SS10[25][33] = 4'hD;
    SS10[26][33] = 4'hD;
    SS10[27][33] = 4'hE;
    SS10[28][33] = 4'hE;
    SS10[29][33] = 4'hE;
    SS10[30][33] = 4'hC;
    SS10[31][33] = 4'hC;
    SS10[32][33] = 4'hC;
    SS10[33][33] = 4'hC;
    SS10[34][33] = 4'hC;
    SS10[35][33] = 4'hC;
    SS10[36][33] = 4'hC;
    SS10[37][33] = 4'hC;
    SS10[38][33] = 4'hC;
    SS10[39][33] = 4'hC;
    SS10[40][33] = 4'hC;
    SS10[41][33] = 4'hC;
    SS10[42][33] = 4'hD;
    SS10[43][33] = 4'hD;
    SS10[44][33] = 4'hD;
    SS10[45][33] = 4'h0;
    SS10[46][33] = 4'h0;
    SS10[47][33] = 4'h0;
    SS10[0][34] = 4'h0;
    SS10[1][34] = 4'h0;
    SS10[2][34] = 4'h0;
    SS10[3][34] = 4'h0;
    SS10[4][34] = 4'h0;
    SS10[5][34] = 4'h0;
    SS10[6][34] = 4'h0;
    SS10[7][34] = 4'h0;
    SS10[8][34] = 4'h0;
    SS10[9][34] = 4'h0;
    SS10[10][34] = 4'h0;
    SS10[11][34] = 4'h0;
    SS10[12][34] = 4'h0;
    SS10[13][34] = 4'h0;
    SS10[14][34] = 4'h0;
    SS10[15][34] = 4'h0;
    SS10[16][34] = 4'h0;
    SS10[17][34] = 4'h0;
    SS10[18][34] = 4'h3;
    SS10[19][34] = 4'h3;
    SS10[20][34] = 4'h3;
    SS10[21][34] = 4'hD;
    SS10[22][34] = 4'hD;
    SS10[23][34] = 4'hD;
    SS10[24][34] = 4'hD;
    SS10[25][34] = 4'hD;
    SS10[26][34] = 4'hD;
    SS10[27][34] = 4'hE;
    SS10[28][34] = 4'hE;
    SS10[29][34] = 4'hE;
    SS10[30][34] = 4'hC;
    SS10[31][34] = 4'hC;
    SS10[32][34] = 4'hC;
    SS10[33][34] = 4'hC;
    SS10[34][34] = 4'hC;
    SS10[35][34] = 4'hC;
    SS10[36][34] = 4'hC;
    SS10[37][34] = 4'hC;
    SS10[38][34] = 4'hC;
    SS10[39][34] = 4'hC;
    SS10[40][34] = 4'hC;
    SS10[41][34] = 4'hC;
    SS10[42][34] = 4'hD;
    SS10[43][34] = 4'hD;
    SS10[44][34] = 4'hD;
    SS10[45][34] = 4'h0;
    SS10[46][34] = 4'h0;
    SS10[47][34] = 4'h0;
    SS10[0][35] = 4'h0;
    SS10[1][35] = 4'h0;
    SS10[2][35] = 4'h0;
    SS10[3][35] = 4'h0;
    SS10[4][35] = 4'h0;
    SS10[5][35] = 4'h0;
    SS10[6][35] = 4'h0;
    SS10[7][35] = 4'h0;
    SS10[8][35] = 4'h0;
    SS10[9][35] = 4'h0;
    SS10[10][35] = 4'h0;
    SS10[11][35] = 4'h0;
    SS10[12][35] = 4'h0;
    SS10[13][35] = 4'h0;
    SS10[14][35] = 4'h0;
    SS10[15][35] = 4'h0;
    SS10[16][35] = 4'h0;
    SS10[17][35] = 4'h0;
    SS10[18][35] = 4'h3;
    SS10[19][35] = 4'h3;
    SS10[20][35] = 4'h3;
    SS10[21][35] = 4'hD;
    SS10[22][35] = 4'hD;
    SS10[23][35] = 4'hD;
    SS10[24][35] = 4'hD;
    SS10[25][35] = 4'hD;
    SS10[26][35] = 4'hD;
    SS10[27][35] = 4'hE;
    SS10[28][35] = 4'hE;
    SS10[29][35] = 4'hE;
    SS10[30][35] = 4'hC;
    SS10[31][35] = 4'hC;
    SS10[32][35] = 4'hC;
    SS10[33][35] = 4'hC;
    SS10[34][35] = 4'hC;
    SS10[35][35] = 4'hC;
    SS10[36][35] = 4'hC;
    SS10[37][35] = 4'hC;
    SS10[38][35] = 4'hC;
    SS10[39][35] = 4'hC;
    SS10[40][35] = 4'hC;
    SS10[41][35] = 4'hC;
    SS10[42][35] = 4'hD;
    SS10[43][35] = 4'hD;
    SS10[44][35] = 4'hD;
    SS10[45][35] = 4'h0;
    SS10[46][35] = 4'h0;
    SS10[47][35] = 4'h0;
    SS10[0][36] = 4'h0;
    SS10[1][36] = 4'h0;
    SS10[2][36] = 4'h0;
    SS10[3][36] = 4'h0;
    SS10[4][36] = 4'h0;
    SS10[5][36] = 4'h0;
    SS10[6][36] = 4'h0;
    SS10[7][36] = 4'h0;
    SS10[8][36] = 4'h0;
    SS10[9][36] = 4'h0;
    SS10[10][36] = 4'h0;
    SS10[11][36] = 4'h0;
    SS10[12][36] = 4'h0;
    SS10[13][36] = 4'h0;
    SS10[14][36] = 4'h0;
    SS10[15][36] = 4'h0;
    SS10[16][36] = 4'h0;
    SS10[17][36] = 4'h0;
    SS10[18][36] = 4'h0;
    SS10[19][36] = 4'h0;
    SS10[20][36] = 4'h0;
    SS10[21][36] = 4'h0;
    SS10[22][36] = 4'h0;
    SS10[23][36] = 4'h0;
    SS10[24][36] = 4'hD;
    SS10[25][36] = 4'hD;
    SS10[26][36] = 4'hD;
    SS10[27][36] = 4'hE;
    SS10[28][36] = 4'hE;
    SS10[29][36] = 4'hE;
    SS10[30][36] = 4'hE;
    SS10[31][36] = 4'hE;
    SS10[32][36] = 4'hE;
    SS10[33][36] = 4'h0;
    SS10[34][36] = 4'h0;
    SS10[35][36] = 4'h0;
    SS10[36][36] = 4'h0;
    SS10[37][36] = 4'h0;
    SS10[38][36] = 4'h0;
    SS10[39][36] = 4'hC;
    SS10[40][36] = 4'hC;
    SS10[41][36] = 4'hC;
    SS10[42][36] = 4'hC;
    SS10[43][36] = 4'hC;
    SS10[44][36] = 4'hC;
    SS10[45][36] = 4'hD;
    SS10[46][36] = 4'hD;
    SS10[47][36] = 4'hD;
    SS10[0][37] = 4'h0;
    SS10[1][37] = 4'h0;
    SS10[2][37] = 4'h0;
    SS10[3][37] = 4'h0;
    SS10[4][37] = 4'h0;
    SS10[5][37] = 4'h0;
    SS10[6][37] = 4'h0;
    SS10[7][37] = 4'h0;
    SS10[8][37] = 4'h0;
    SS10[9][37] = 4'h0;
    SS10[10][37] = 4'h0;
    SS10[11][37] = 4'h0;
    SS10[12][37] = 4'h0;
    SS10[13][37] = 4'h0;
    SS10[14][37] = 4'h0;
    SS10[15][37] = 4'h0;
    SS10[16][37] = 4'h0;
    SS10[17][37] = 4'h0;
    SS10[18][37] = 4'h0;
    SS10[19][37] = 4'h0;
    SS10[20][37] = 4'h0;
    SS10[21][37] = 4'h0;
    SS10[22][37] = 4'h0;
    SS10[23][37] = 4'h0;
    SS10[24][37] = 4'hD;
    SS10[25][37] = 4'hD;
    SS10[26][37] = 4'hD;
    SS10[27][37] = 4'hE;
    SS10[28][37] = 4'hE;
    SS10[29][37] = 4'hE;
    SS10[30][37] = 4'hE;
    SS10[31][37] = 4'hE;
    SS10[32][37] = 4'hE;
    SS10[33][37] = 4'h0;
    SS10[34][37] = 4'h0;
    SS10[35][37] = 4'h0;
    SS10[36][37] = 4'h0;
    SS10[37][37] = 4'h0;
    SS10[38][37] = 4'h0;
    SS10[39][37] = 4'hC;
    SS10[40][37] = 4'hC;
    SS10[41][37] = 4'hC;
    SS10[42][37] = 4'hC;
    SS10[43][37] = 4'hC;
    SS10[44][37] = 4'hC;
    SS10[45][37] = 4'hD;
    SS10[46][37] = 4'hD;
    SS10[47][37] = 4'hD;
    SS10[0][38] = 4'h0;
    SS10[1][38] = 4'h0;
    SS10[2][38] = 4'h0;
    SS10[3][38] = 4'h0;
    SS10[4][38] = 4'h0;
    SS10[5][38] = 4'h0;
    SS10[6][38] = 4'h0;
    SS10[7][38] = 4'h0;
    SS10[8][38] = 4'h0;
    SS10[9][38] = 4'h0;
    SS10[10][38] = 4'h0;
    SS10[11][38] = 4'h0;
    SS10[12][38] = 4'h0;
    SS10[13][38] = 4'h0;
    SS10[14][38] = 4'h0;
    SS10[15][38] = 4'h0;
    SS10[16][38] = 4'h0;
    SS10[17][38] = 4'h0;
    SS10[18][38] = 4'h0;
    SS10[19][38] = 4'h0;
    SS10[20][38] = 4'h0;
    SS10[21][38] = 4'h0;
    SS10[22][38] = 4'h0;
    SS10[23][38] = 4'h0;
    SS10[24][38] = 4'hD;
    SS10[25][38] = 4'hD;
    SS10[26][38] = 4'hD;
    SS10[27][38] = 4'hE;
    SS10[28][38] = 4'hE;
    SS10[29][38] = 4'hE;
    SS10[30][38] = 4'hE;
    SS10[31][38] = 4'hE;
    SS10[32][38] = 4'hE;
    SS10[33][38] = 4'h0;
    SS10[34][38] = 4'h0;
    SS10[35][38] = 4'h0;
    SS10[36][38] = 4'h0;
    SS10[37][38] = 4'h0;
    SS10[38][38] = 4'h0;
    SS10[39][38] = 4'hC;
    SS10[40][38] = 4'hC;
    SS10[41][38] = 4'hC;
    SS10[42][38] = 4'hC;
    SS10[43][38] = 4'hC;
    SS10[44][38] = 4'hC;
    SS10[45][38] = 4'hD;
    SS10[46][38] = 4'hD;
    SS10[47][38] = 4'hD;
    SS10[0][39] = 4'h0;
    SS10[1][39] = 4'h0;
    SS10[2][39] = 4'h0;
    SS10[3][39] = 4'h0;
    SS10[4][39] = 4'h0;
    SS10[5][39] = 4'h0;
    SS10[6][39] = 4'h0;
    SS10[7][39] = 4'h0;
    SS10[8][39] = 4'h0;
    SS10[9][39] = 4'h0;
    SS10[10][39] = 4'h0;
    SS10[11][39] = 4'h0;
    SS10[12][39] = 4'h0;
    SS10[13][39] = 4'h0;
    SS10[14][39] = 4'h0;
    SS10[15][39] = 4'h0;
    SS10[16][39] = 4'h0;
    SS10[17][39] = 4'h0;
    SS10[18][39] = 4'h0;
    SS10[19][39] = 4'h0;
    SS10[20][39] = 4'h0;
    SS10[21][39] = 4'h0;
    SS10[22][39] = 4'h0;
    SS10[23][39] = 4'h0;
    SS10[24][39] = 4'h3;
    SS10[25][39] = 4'h3;
    SS10[26][39] = 4'h3;
    SS10[27][39] = 4'hD;
    SS10[28][39] = 4'hD;
    SS10[29][39] = 4'hD;
    SS10[30][39] = 4'hE;
    SS10[31][39] = 4'hE;
    SS10[32][39] = 4'hE;
    SS10[33][39] = 4'h0;
    SS10[34][39] = 4'h0;
    SS10[35][39] = 4'h0;
    SS10[36][39] = 4'h0;
    SS10[37][39] = 4'h0;
    SS10[38][39] = 4'h0;
    SS10[39][39] = 4'h0;
    SS10[40][39] = 4'h0;
    SS10[41][39] = 4'h0;
    SS10[42][39] = 4'h0;
    SS10[43][39] = 4'h0;
    SS10[44][39] = 4'h0;
    SS10[45][39] = 4'h0;
    SS10[46][39] = 4'h0;
    SS10[47][39] = 4'h0;
    SS10[0][40] = 4'h0;
    SS10[1][40] = 4'h0;
    SS10[2][40] = 4'h0;
    SS10[3][40] = 4'h0;
    SS10[4][40] = 4'h0;
    SS10[5][40] = 4'h0;
    SS10[6][40] = 4'h0;
    SS10[7][40] = 4'h0;
    SS10[8][40] = 4'h0;
    SS10[9][40] = 4'h0;
    SS10[10][40] = 4'h0;
    SS10[11][40] = 4'h0;
    SS10[12][40] = 4'h0;
    SS10[13][40] = 4'h0;
    SS10[14][40] = 4'h0;
    SS10[15][40] = 4'h0;
    SS10[16][40] = 4'h0;
    SS10[17][40] = 4'h0;
    SS10[18][40] = 4'h0;
    SS10[19][40] = 4'h0;
    SS10[20][40] = 4'h0;
    SS10[21][40] = 4'h0;
    SS10[22][40] = 4'h0;
    SS10[23][40] = 4'h0;
    SS10[24][40] = 4'h3;
    SS10[25][40] = 4'h3;
    SS10[26][40] = 4'h3;
    SS10[27][40] = 4'hD;
    SS10[28][40] = 4'hD;
    SS10[29][40] = 4'hD;
    SS10[30][40] = 4'hE;
    SS10[31][40] = 4'hE;
    SS10[32][40] = 4'hE;
    SS10[33][40] = 4'h0;
    SS10[34][40] = 4'h0;
    SS10[35][40] = 4'h0;
    SS10[36][40] = 4'h0;
    SS10[37][40] = 4'h0;
    SS10[38][40] = 4'h0;
    SS10[39][40] = 4'h0;
    SS10[40][40] = 4'h0;
    SS10[41][40] = 4'h0;
    SS10[42][40] = 4'h0;
    SS10[43][40] = 4'h0;
    SS10[44][40] = 4'h0;
    SS10[45][40] = 4'h0;
    SS10[46][40] = 4'h0;
    SS10[47][40] = 4'h0;
    SS10[0][41] = 4'h0;
    SS10[1][41] = 4'h0;
    SS10[2][41] = 4'h0;
    SS10[3][41] = 4'h0;
    SS10[4][41] = 4'h0;
    SS10[5][41] = 4'h0;
    SS10[6][41] = 4'h0;
    SS10[7][41] = 4'h0;
    SS10[8][41] = 4'h0;
    SS10[9][41] = 4'h0;
    SS10[10][41] = 4'h0;
    SS10[11][41] = 4'h0;
    SS10[12][41] = 4'h0;
    SS10[13][41] = 4'h0;
    SS10[14][41] = 4'h0;
    SS10[15][41] = 4'h0;
    SS10[16][41] = 4'h0;
    SS10[17][41] = 4'h0;
    SS10[18][41] = 4'h0;
    SS10[19][41] = 4'h0;
    SS10[20][41] = 4'h0;
    SS10[21][41] = 4'h0;
    SS10[22][41] = 4'h0;
    SS10[23][41] = 4'h0;
    SS10[24][41] = 4'h3;
    SS10[25][41] = 4'h3;
    SS10[26][41] = 4'h3;
    SS10[27][41] = 4'hD;
    SS10[28][41] = 4'hD;
    SS10[29][41] = 4'hD;
    SS10[30][41] = 4'hE;
    SS10[31][41] = 4'hE;
    SS10[32][41] = 4'hE;
    SS10[33][41] = 4'h0;
    SS10[34][41] = 4'h0;
    SS10[35][41] = 4'h0;
    SS10[36][41] = 4'h0;
    SS10[37][41] = 4'h0;
    SS10[38][41] = 4'h0;
    SS10[39][41] = 4'h0;
    SS10[40][41] = 4'h0;
    SS10[41][41] = 4'h0;
    SS10[42][41] = 4'h0;
    SS10[43][41] = 4'h0;
    SS10[44][41] = 4'h0;
    SS10[45][41] = 4'h0;
    SS10[46][41] = 4'h0;
    SS10[47][41] = 4'h0;
    SS10[0][42] = 4'h0;
    SS10[1][42] = 4'h0;
    SS10[2][42] = 4'h0;
    SS10[3][42] = 4'h0;
    SS10[4][42] = 4'h0;
    SS10[5][42] = 4'h0;
    SS10[6][42] = 4'h0;
    SS10[7][42] = 4'h0;
    SS10[8][42] = 4'h0;
    SS10[9][42] = 4'h0;
    SS10[10][42] = 4'h0;
    SS10[11][42] = 4'h0;
    SS10[12][42] = 4'h0;
    SS10[13][42] = 4'h0;
    SS10[14][42] = 4'h0;
    SS10[15][42] = 4'h0;
    SS10[16][42] = 4'h0;
    SS10[17][42] = 4'h0;
    SS10[18][42] = 4'h0;
    SS10[19][42] = 4'h0;
    SS10[20][42] = 4'h0;
    SS10[21][42] = 4'h0;
    SS10[22][42] = 4'h0;
    SS10[23][42] = 4'h0;
    SS10[24][42] = 4'h0;
    SS10[25][42] = 4'h0;
    SS10[26][42] = 4'h0;
    SS10[27][42] = 4'hD;
    SS10[28][42] = 4'hD;
    SS10[29][42] = 4'hD;
    SS10[30][42] = 4'hD;
    SS10[31][42] = 4'hD;
    SS10[32][42] = 4'hD;
    SS10[33][42] = 4'h0;
    SS10[34][42] = 4'h0;
    SS10[35][42] = 4'h0;
    SS10[36][42] = 4'h0;
    SS10[37][42] = 4'h0;
    SS10[38][42] = 4'h0;
    SS10[39][42] = 4'h0;
    SS10[40][42] = 4'h0;
    SS10[41][42] = 4'h0;
    SS10[42][42] = 4'h0;
    SS10[43][42] = 4'h0;
    SS10[44][42] = 4'h0;
    SS10[45][42] = 4'h0;
    SS10[46][42] = 4'h0;
    SS10[47][42] = 4'h0;
    SS10[0][43] = 4'h0;
    SS10[1][43] = 4'h0;
    SS10[2][43] = 4'h0;
    SS10[3][43] = 4'h0;
    SS10[4][43] = 4'h0;
    SS10[5][43] = 4'h0;
    SS10[6][43] = 4'h0;
    SS10[7][43] = 4'h0;
    SS10[8][43] = 4'h0;
    SS10[9][43] = 4'h0;
    SS10[10][43] = 4'h0;
    SS10[11][43] = 4'h0;
    SS10[12][43] = 4'h0;
    SS10[13][43] = 4'h0;
    SS10[14][43] = 4'h0;
    SS10[15][43] = 4'h0;
    SS10[16][43] = 4'h0;
    SS10[17][43] = 4'h0;
    SS10[18][43] = 4'h0;
    SS10[19][43] = 4'h0;
    SS10[20][43] = 4'h0;
    SS10[21][43] = 4'h0;
    SS10[22][43] = 4'h0;
    SS10[23][43] = 4'h0;
    SS10[24][43] = 4'h0;
    SS10[25][43] = 4'h0;
    SS10[26][43] = 4'h0;
    SS10[27][43] = 4'hD;
    SS10[28][43] = 4'hD;
    SS10[29][43] = 4'hD;
    SS10[30][43] = 4'hD;
    SS10[31][43] = 4'hD;
    SS10[32][43] = 4'hD;
    SS10[33][43] = 4'h0;
    SS10[34][43] = 4'h0;
    SS10[35][43] = 4'h0;
    SS10[36][43] = 4'h0;
    SS10[37][43] = 4'h0;
    SS10[38][43] = 4'h0;
    SS10[39][43] = 4'h0;
    SS10[40][43] = 4'h0;
    SS10[41][43] = 4'h0;
    SS10[42][43] = 4'h0;
    SS10[43][43] = 4'h0;
    SS10[44][43] = 4'h0;
    SS10[45][43] = 4'h0;
    SS10[46][43] = 4'h0;
    SS10[47][43] = 4'h0;
    SS10[0][44] = 4'h0;
    SS10[1][44] = 4'h0;
    SS10[2][44] = 4'h0;
    SS10[3][44] = 4'h0;
    SS10[4][44] = 4'h0;
    SS10[5][44] = 4'h0;
    SS10[6][44] = 4'h0;
    SS10[7][44] = 4'h0;
    SS10[8][44] = 4'h0;
    SS10[9][44] = 4'h0;
    SS10[10][44] = 4'h0;
    SS10[11][44] = 4'h0;
    SS10[12][44] = 4'h0;
    SS10[13][44] = 4'h0;
    SS10[14][44] = 4'h0;
    SS10[15][44] = 4'h0;
    SS10[16][44] = 4'h0;
    SS10[17][44] = 4'h0;
    SS10[18][44] = 4'h0;
    SS10[19][44] = 4'h0;
    SS10[20][44] = 4'h0;
    SS10[21][44] = 4'h0;
    SS10[22][44] = 4'h0;
    SS10[23][44] = 4'h0;
    SS10[24][44] = 4'h0;
    SS10[25][44] = 4'h0;
    SS10[26][44] = 4'h0;
    SS10[27][44] = 4'hD;
    SS10[28][44] = 4'hD;
    SS10[29][44] = 4'hD;
    SS10[30][44] = 4'hD;
    SS10[31][44] = 4'hD;
    SS10[32][44] = 4'hD;
    SS10[33][44] = 4'h0;
    SS10[34][44] = 4'h0;
    SS10[35][44] = 4'h0;
    SS10[36][44] = 4'h0;
    SS10[37][44] = 4'h0;
    SS10[38][44] = 4'h0;
    SS10[39][44] = 4'h0;
    SS10[40][44] = 4'h0;
    SS10[41][44] = 4'h0;
    SS10[42][44] = 4'h0;
    SS10[43][44] = 4'h0;
    SS10[44][44] = 4'h0;
    SS10[45][44] = 4'h0;
    SS10[46][44] = 4'h0;
    SS10[47][44] = 4'h0;
    SS10[0][45] = 4'h0;
    SS10[1][45] = 4'h0;
    SS10[2][45] = 4'h0;
    SS10[3][45] = 4'h0;
    SS10[4][45] = 4'h0;
    SS10[5][45] = 4'h0;
    SS10[6][45] = 4'h0;
    SS10[7][45] = 4'h0;
    SS10[8][45] = 4'h0;
    SS10[9][45] = 4'h0;
    SS10[10][45] = 4'h0;
    SS10[11][45] = 4'h0;
    SS10[12][45] = 4'h0;
    SS10[13][45] = 4'h0;
    SS10[14][45] = 4'h0;
    SS10[15][45] = 4'h0;
    SS10[16][45] = 4'h0;
    SS10[17][45] = 4'h0;
    SS10[18][45] = 4'h0;
    SS10[19][45] = 4'h0;
    SS10[20][45] = 4'h0;
    SS10[21][45] = 4'h0;
    SS10[22][45] = 4'h0;
    SS10[23][45] = 4'h0;
    SS10[24][45] = 4'h0;
    SS10[25][45] = 4'h0;
    SS10[26][45] = 4'h0;
    SS10[27][45] = 4'h0;
    SS10[28][45] = 4'h0;
    SS10[29][45] = 4'h0;
    SS10[30][45] = 4'hD;
    SS10[31][45] = 4'hD;
    SS10[32][45] = 4'hD;
    SS10[33][45] = 4'h0;
    SS10[34][45] = 4'h0;
    SS10[35][45] = 4'h0;
    SS10[36][45] = 4'h0;
    SS10[37][45] = 4'h0;
    SS10[38][45] = 4'h0;
    SS10[39][45] = 4'h0;
    SS10[40][45] = 4'h0;
    SS10[41][45] = 4'h0;
    SS10[42][45] = 4'h0;
    SS10[43][45] = 4'h0;
    SS10[44][45] = 4'h0;
    SS10[45][45] = 4'h0;
    SS10[46][45] = 4'h0;
    SS10[47][45] = 4'h0;
    SS10[0][46] = 4'h0;
    SS10[1][46] = 4'h0;
    SS10[2][46] = 4'h0;
    SS10[3][46] = 4'h0;
    SS10[4][46] = 4'h0;
    SS10[5][46] = 4'h0;
    SS10[6][46] = 4'h0;
    SS10[7][46] = 4'h0;
    SS10[8][46] = 4'h0;
    SS10[9][46] = 4'h0;
    SS10[10][46] = 4'h0;
    SS10[11][46] = 4'h0;
    SS10[12][46] = 4'h0;
    SS10[13][46] = 4'h0;
    SS10[14][46] = 4'h0;
    SS10[15][46] = 4'h0;
    SS10[16][46] = 4'h0;
    SS10[17][46] = 4'h0;
    SS10[18][46] = 4'h0;
    SS10[19][46] = 4'h0;
    SS10[20][46] = 4'h0;
    SS10[21][46] = 4'h0;
    SS10[22][46] = 4'h0;
    SS10[23][46] = 4'h0;
    SS10[24][46] = 4'h0;
    SS10[25][46] = 4'h0;
    SS10[26][46] = 4'h0;
    SS10[27][46] = 4'h0;
    SS10[28][46] = 4'h0;
    SS10[29][46] = 4'h0;
    SS10[30][46] = 4'hD;
    SS10[31][46] = 4'hD;
    SS10[32][46] = 4'hD;
    SS10[33][46] = 4'h0;
    SS10[34][46] = 4'h0;
    SS10[35][46] = 4'h0;
    SS10[36][46] = 4'h0;
    SS10[37][46] = 4'h0;
    SS10[38][46] = 4'h0;
    SS10[39][46] = 4'h0;
    SS10[40][46] = 4'h0;
    SS10[41][46] = 4'h0;
    SS10[42][46] = 4'h0;
    SS10[43][46] = 4'h0;
    SS10[44][46] = 4'h0;
    SS10[45][46] = 4'h0;
    SS10[46][46] = 4'h0;
    SS10[47][46] = 4'h0;
    SS10[0][47] = 4'h0;
    SS10[1][47] = 4'h0;
    SS10[2][47] = 4'h0;
    SS10[3][47] = 4'h0;
    SS10[4][47] = 4'h0;
    SS10[5][47] = 4'h0;
    SS10[6][47] = 4'h0;
    SS10[7][47] = 4'h0;
    SS10[8][47] = 4'h0;
    SS10[9][47] = 4'h0;
    SS10[10][47] = 4'h0;
    SS10[11][47] = 4'h0;
    SS10[12][47] = 4'h0;
    SS10[13][47] = 4'h0;
    SS10[14][47] = 4'h0;
    SS10[15][47] = 4'h0;
    SS10[16][47] = 4'h0;
    SS10[17][47] = 4'h0;
    SS10[18][47] = 4'h0;
    SS10[19][47] = 4'h0;
    SS10[20][47] = 4'h0;
    SS10[21][47] = 4'h0;
    SS10[22][47] = 4'h0;
    SS10[23][47] = 4'h0;
    SS10[24][47] = 4'h0;
    SS10[25][47] = 4'h0;
    SS10[26][47] = 4'h0;
    SS10[27][47] = 4'h0;
    SS10[28][47] = 4'h0;
    SS10[29][47] = 4'h0;
    SS10[30][47] = 4'hD;
    SS10[31][47] = 4'hD;
    SS10[32][47] = 4'hD;
    SS10[33][47] = 4'h0;
    SS10[34][47] = 4'h0;
    SS10[35][47] = 4'h0;
    SS10[36][47] = 4'h0;
    SS10[37][47] = 4'h0;
    SS10[38][47] = 4'h0;
    SS10[39][47] = 4'h0;
    SS10[40][47] = 4'h0;
    SS10[41][47] = 4'h0;
    SS10[42][47] = 4'h0;
    SS10[43][47] = 4'h0;
    SS10[44][47] = 4'h0;
    SS10[45][47] = 4'h0;
    SS10[46][47] = 4'h0;
    SS10[47][47] = 4'h0;
 
//SS 11
    SS11[0][0] = 4'h0;
    SS11[1][0] = 4'h0;
    SS11[2][0] = 4'h0;
    SS11[3][0] = 4'h0;
    SS11[4][0] = 4'h0;
    SS11[5][0] = 4'h0;
    SS11[6][0] = 4'h0;
    SS11[7][0] = 4'h0;
    SS11[8][0] = 4'h0;
    SS11[9][0] = 4'h0;
    SS11[10][0] = 4'h0;
    SS11[11][0] = 4'h0;
    SS11[12][0] = 4'h0;
    SS11[13][0] = 4'h0;
    SS11[14][0] = 4'h0;
    SS11[15][0] = 4'h0;
    SS11[16][0] = 4'h0;
    SS11[17][0] = 4'h0;
    SS11[18][0] = 4'h0;
    SS11[19][0] = 4'h0;
    SS11[20][0] = 4'h0;
    SS11[21][0] = 4'h0;
    SS11[22][0] = 4'h0;
    SS11[23][0] = 4'h0;
    SS11[24][0] = 4'h0;
    SS11[25][0] = 4'h0;
    SS11[26][0] = 4'h0;
    SS11[27][0] = 4'h0;
    SS11[28][0] = 4'h0;
    SS11[29][0] = 4'h0;
    SS11[30][0] = 4'h0;
    SS11[31][0] = 4'h0;
    SS11[32][0] = 4'h0;
    SS11[33][0] = 4'h0;
    SS11[34][0] = 4'h0;
    SS11[35][0] = 4'h0;
    SS11[36][0] = 4'h0;
    SS11[37][0] = 4'h0;
    SS11[38][0] = 4'h0;
    SS11[39][0] = 4'h0;
    SS11[40][0] = 4'h0;
    SS11[41][0] = 4'h0;
    SS11[42][0] = 4'h0;
    SS11[43][0] = 4'h0;
    SS11[44][0] = 4'h0;
    SS11[45][0] = 4'h0;
    SS11[46][0] = 4'h0;
    SS11[47][0] = 4'h0;
    SS11[0][1] = 4'h0;
    SS11[1][1] = 4'h0;
    SS11[2][1] = 4'h0;
    SS11[3][1] = 4'h0;
    SS11[4][1] = 4'h0;
    SS11[5][1] = 4'h0;
    SS11[6][1] = 4'h0;
    SS11[7][1] = 4'h0;
    SS11[8][1] = 4'h0;
    SS11[9][1] = 4'h0;
    SS11[10][1] = 4'h0;
    SS11[11][1] = 4'h0;
    SS11[12][1] = 4'h0;
    SS11[13][1] = 4'h0;
    SS11[14][1] = 4'h0;
    SS11[15][1] = 4'h0;
    SS11[16][1] = 4'h0;
    SS11[17][1] = 4'h0;
    SS11[18][1] = 4'h0;
    SS11[19][1] = 4'h0;
    SS11[20][1] = 4'h0;
    SS11[21][1] = 4'h0;
    SS11[22][1] = 4'h0;
    SS11[23][1] = 4'h0;
    SS11[24][1] = 4'h0;
    SS11[25][1] = 4'h0;
    SS11[26][1] = 4'h0;
    SS11[27][1] = 4'h0;
    SS11[28][1] = 4'h0;
    SS11[29][1] = 4'h0;
    SS11[30][1] = 4'h0;
    SS11[31][1] = 4'h0;
    SS11[32][1] = 4'h0;
    SS11[33][1] = 4'h0;
    SS11[34][1] = 4'h0;
    SS11[35][1] = 4'h0;
    SS11[36][1] = 4'h0;
    SS11[37][1] = 4'h0;
    SS11[38][1] = 4'h0;
    SS11[39][1] = 4'h0;
    SS11[40][1] = 4'h0;
    SS11[41][1] = 4'h0;
    SS11[42][1] = 4'h0;
    SS11[43][1] = 4'h0;
    SS11[44][1] = 4'h0;
    SS11[45][1] = 4'h0;
    SS11[46][1] = 4'h0;
    SS11[47][1] = 4'h0;
    SS11[0][2] = 4'h0;
    SS11[1][2] = 4'h0;
    SS11[2][2] = 4'h0;
    SS11[3][2] = 4'h0;
    SS11[4][2] = 4'h0;
    SS11[5][2] = 4'h0;
    SS11[6][2] = 4'h0;
    SS11[7][2] = 4'h0;
    SS11[8][2] = 4'h0;
    SS11[9][2] = 4'h0;
    SS11[10][2] = 4'h0;
    SS11[11][2] = 4'h0;
    SS11[12][2] = 4'h0;
    SS11[13][2] = 4'h0;
    SS11[14][2] = 4'h0;
    SS11[15][2] = 4'h0;
    SS11[16][2] = 4'h0;
    SS11[17][2] = 4'h0;
    SS11[18][2] = 4'h0;
    SS11[19][2] = 4'h0;
    SS11[20][2] = 4'h0;
    SS11[21][2] = 4'h0;
    SS11[22][2] = 4'h0;
    SS11[23][2] = 4'h0;
    SS11[24][2] = 4'h0;
    SS11[25][2] = 4'h0;
    SS11[26][2] = 4'h0;
    SS11[27][2] = 4'h0;
    SS11[28][2] = 4'h0;
    SS11[29][2] = 4'h0;
    SS11[30][2] = 4'h0;
    SS11[31][2] = 4'h0;
    SS11[32][2] = 4'h0;
    SS11[33][2] = 4'h0;
    SS11[34][2] = 4'h0;
    SS11[35][2] = 4'h0;
    SS11[36][2] = 4'h0;
    SS11[37][2] = 4'h0;
    SS11[38][2] = 4'h0;
    SS11[39][2] = 4'h0;
    SS11[40][2] = 4'h0;
    SS11[41][2] = 4'h0;
    SS11[42][2] = 4'h0;
    SS11[43][2] = 4'h0;
    SS11[44][2] = 4'h0;
    SS11[45][2] = 4'h0;
    SS11[46][2] = 4'h0;
    SS11[47][2] = 4'h0;
    SS11[0][3] = 4'h0;
    SS11[1][3] = 4'h0;
    SS11[2][3] = 4'h0;
    SS11[3][3] = 4'h0;
    SS11[4][3] = 4'h0;
    SS11[5][3] = 4'h0;
    SS11[6][3] = 4'h0;
    SS11[7][3] = 4'h0;
    SS11[8][3] = 4'h0;
    SS11[9][3] = 4'h0;
    SS11[10][3] = 4'h0;
    SS11[11][3] = 4'h0;
    SS11[12][3] = 4'h0;
    SS11[13][3] = 4'h0;
    SS11[14][3] = 4'h0;
    SS11[15][3] = 4'h0;
    SS11[16][3] = 4'h0;
    SS11[17][3] = 4'h0;
    SS11[18][3] = 4'h0;
    SS11[19][3] = 4'h0;
    SS11[20][3] = 4'h0;
    SS11[21][3] = 4'h0;
    SS11[22][3] = 4'h0;
    SS11[23][3] = 4'h0;
    SS11[24][3] = 4'h0;
    SS11[25][3] = 4'h0;
    SS11[26][3] = 4'h0;
    SS11[27][3] = 4'h0;
    SS11[28][3] = 4'h0;
    SS11[29][3] = 4'h0;
    SS11[30][3] = 4'h0;
    SS11[31][3] = 4'h0;
    SS11[32][3] = 4'h0;
    SS11[33][3] = 4'h0;
    SS11[34][3] = 4'h0;
    SS11[35][3] = 4'h0;
    SS11[36][3] = 4'h0;
    SS11[37][3] = 4'h0;
    SS11[38][3] = 4'h0;
    SS11[39][3] = 4'h0;
    SS11[40][3] = 4'h0;
    SS11[41][3] = 4'h0;
    SS11[42][3] = 4'h0;
    SS11[43][3] = 4'h0;
    SS11[44][3] = 4'h0;
    SS11[45][3] = 4'h0;
    SS11[46][3] = 4'h0;
    SS11[47][3] = 4'h0;
    SS11[0][4] = 4'h0;
    SS11[1][4] = 4'h0;
    SS11[2][4] = 4'h0;
    SS11[3][4] = 4'h0;
    SS11[4][4] = 4'h0;
    SS11[5][4] = 4'h0;
    SS11[6][4] = 4'h0;
    SS11[7][4] = 4'h0;
    SS11[8][4] = 4'h0;
    SS11[9][4] = 4'h0;
    SS11[10][4] = 4'h0;
    SS11[11][4] = 4'h0;
    SS11[12][4] = 4'h0;
    SS11[13][4] = 4'h0;
    SS11[14][4] = 4'h0;
    SS11[15][4] = 4'h0;
    SS11[16][4] = 4'h0;
    SS11[17][4] = 4'h0;
    SS11[18][4] = 4'h0;
    SS11[19][4] = 4'h0;
    SS11[20][4] = 4'h0;
    SS11[21][4] = 4'h0;
    SS11[22][4] = 4'h0;
    SS11[23][4] = 4'h0;
    SS11[24][4] = 4'h0;
    SS11[25][4] = 4'h0;
    SS11[26][4] = 4'h0;
    SS11[27][4] = 4'h0;
    SS11[28][4] = 4'h0;
    SS11[29][4] = 4'h0;
    SS11[30][4] = 4'h0;
    SS11[31][4] = 4'h0;
    SS11[32][4] = 4'h0;
    SS11[33][4] = 4'h0;
    SS11[34][4] = 4'h0;
    SS11[35][4] = 4'h0;
    SS11[36][4] = 4'h0;
    SS11[37][4] = 4'h0;
    SS11[38][4] = 4'hD;
    SS11[39][4] = 4'h0;
    SS11[40][4] = 4'h0;
    SS11[41][4] = 4'h0;
    SS11[42][4] = 4'h0;
    SS11[43][4] = 4'h0;
    SS11[44][4] = 4'h0;
    SS11[45][4] = 4'h0;
    SS11[46][4] = 4'h0;
    SS11[47][4] = 4'h0;
    SS11[0][5] = 4'h0;
    SS11[1][5] = 4'h0;
    SS11[2][5] = 4'h0;
    SS11[3][5] = 4'h0;
    SS11[4][5] = 4'h0;
    SS11[5][5] = 4'h0;
    SS11[6][5] = 4'h0;
    SS11[7][5] = 4'h0;
    SS11[8][5] = 4'h0;
    SS11[9][5] = 4'h0;
    SS11[10][5] = 4'h0;
    SS11[11][5] = 4'h0;
    SS11[12][5] = 4'h0;
    SS11[13][5] = 4'h0;
    SS11[14][5] = 4'h0;
    SS11[15][5] = 4'h0;
    SS11[16][5] = 4'h0;
    SS11[17][5] = 4'h0;
    SS11[18][5] = 4'h0;
    SS11[19][5] = 4'h0;
    SS11[20][5] = 4'h0;
    SS11[21][5] = 4'h0;
    SS11[22][5] = 4'h0;
    SS11[23][5] = 4'h0;
    SS11[24][5] = 4'h0;
    SS11[25][5] = 4'h0;
    SS11[26][5] = 4'h0;
    SS11[27][5] = 4'h0;
    SS11[28][5] = 4'h0;
    SS11[29][5] = 4'h0;
    SS11[30][5] = 4'h0;
    SS11[31][5] = 4'h0;
    SS11[32][5] = 4'h0;
    SS11[33][5] = 4'h0;
    SS11[34][5] = 4'h0;
    SS11[35][5] = 4'h0;
    SS11[36][5] = 4'h0;
    SS11[37][5] = 4'h0;
    SS11[38][5] = 4'hD;
    SS11[39][5] = 4'hD;
    SS11[40][5] = 4'hD;
    SS11[41][5] = 4'h0;
    SS11[42][5] = 4'h0;
    SS11[43][5] = 4'h0;
    SS11[44][5] = 4'h0;
    SS11[45][5] = 4'h0;
    SS11[46][5] = 4'h0;
    SS11[47][5] = 4'h0;
    SS11[0][6] = 4'h0;
    SS11[1][6] = 4'h0;
    SS11[2][6] = 4'h0;
    SS11[3][6] = 4'h0;
    SS11[4][6] = 4'h0;
    SS11[5][6] = 4'h0;
    SS11[6][6] = 4'h0;
    SS11[7][6] = 4'h0;
    SS11[8][6] = 4'h0;
    SS11[9][6] = 4'h0;
    SS11[10][6] = 4'h0;
    SS11[11][6] = 4'h0;
    SS11[12][6] = 4'h0;
    SS11[13][6] = 4'h0;
    SS11[14][6] = 4'h0;
    SS11[15][6] = 4'h0;
    SS11[16][6] = 4'h0;
    SS11[17][6] = 4'h0;
    SS11[18][6] = 4'h0;
    SS11[19][6] = 4'h0;
    SS11[20][6] = 4'h0;
    SS11[21][6] = 4'h0;
    SS11[22][6] = 4'h0;
    SS11[23][6] = 4'h0;
    SS11[24][6] = 4'h0;
    SS11[25][6] = 4'h0;
    SS11[26][6] = 4'h0;
    SS11[27][6] = 4'h0;
    SS11[28][6] = 4'h0;
    SS11[29][6] = 4'h0;
    SS11[30][6] = 4'h0;
    SS11[31][6] = 4'h0;
    SS11[32][6] = 4'h0;
    SS11[33][6] = 4'h0;
    SS11[34][6] = 4'hD;
    SS11[35][6] = 4'hD;
    SS11[36][6] = 4'h0;
    SS11[37][6] = 4'h0;
    SS11[38][6] = 4'hD;
    SS11[39][6] = 4'hD;
    SS11[40][6] = 4'hD;
    SS11[41][6] = 4'h0;
    SS11[42][6] = 4'h0;
    SS11[43][6] = 4'h0;
    SS11[44][6] = 4'h0;
    SS11[45][6] = 4'h0;
    SS11[46][6] = 4'h0;
    SS11[47][6] = 4'h0;
    SS11[0][7] = 4'h0;
    SS11[1][7] = 4'h0;
    SS11[2][7] = 4'h0;
    SS11[3][7] = 4'h0;
    SS11[4][7] = 4'h0;
    SS11[5][7] = 4'h0;
    SS11[6][7] = 4'h0;
    SS11[7][7] = 4'h0;
    SS11[8][7] = 4'h0;
    SS11[9][7] = 4'h0;
    SS11[10][7] = 4'h0;
    SS11[11][7] = 4'h0;
    SS11[12][7] = 4'h0;
    SS11[13][7] = 4'h0;
    SS11[14][7] = 4'h0;
    SS11[15][7] = 4'h0;
    SS11[16][7] = 4'h0;
    SS11[17][7] = 4'h0;
    SS11[18][7] = 4'h0;
    SS11[19][7] = 4'h0;
    SS11[20][7] = 4'h0;
    SS11[21][7] = 4'h0;
    SS11[22][7] = 4'h0;
    SS11[23][7] = 4'h0;
    SS11[24][7] = 4'h0;
    SS11[25][7] = 4'h0;
    SS11[26][7] = 4'h0;
    SS11[27][7] = 4'h0;
    SS11[28][7] = 4'h0;
    SS11[29][7] = 4'h0;
    SS11[30][7] = 4'h0;
    SS11[31][7] = 4'h0;
    SS11[32][7] = 4'h0;
    SS11[33][7] = 4'h0;
    SS11[34][7] = 4'hD;
    SS11[35][7] = 4'hD;
    SS11[36][7] = 4'hD;
    SS11[37][7] = 4'hD;
    SS11[38][7] = 4'hD;
    SS11[39][7] = 4'hD;
    SS11[40][7] = 4'h0;
    SS11[41][7] = 4'h0;
    SS11[42][7] = 4'h0;
    SS11[43][7] = 4'h0;
    SS11[44][7] = 4'h0;
    SS11[45][7] = 4'h0;
    SS11[46][7] = 4'h0;
    SS11[47][7] = 4'h0;
    SS11[0][8] = 4'h0;
    SS11[1][8] = 4'h0;
    SS11[2][8] = 4'h0;
    SS11[3][8] = 4'h0;
    SS11[4][8] = 4'h0;
    SS11[5][8] = 4'h0;
    SS11[6][8] = 4'h0;
    SS11[7][8] = 4'h0;
    SS11[8][8] = 4'h0;
    SS11[9][8] = 4'h0;
    SS11[10][8] = 4'h0;
    SS11[11][8] = 4'h0;
    SS11[12][8] = 4'h0;
    SS11[13][8] = 4'h0;
    SS11[14][8] = 4'h0;
    SS11[15][8] = 4'h0;
    SS11[16][8] = 4'h0;
    SS11[17][8] = 4'h0;
    SS11[18][8] = 4'h0;
    SS11[19][8] = 4'h0;
    SS11[20][8] = 4'h0;
    SS11[21][8] = 4'h0;
    SS11[22][8] = 4'h0;
    SS11[23][8] = 4'h0;
    SS11[24][8] = 4'h0;
    SS11[25][8] = 4'h0;
    SS11[26][8] = 4'h0;
    SS11[27][8] = 4'h0;
    SS11[28][8] = 4'h0;
    SS11[29][8] = 4'h0;
    SS11[30][8] = 4'h3;
    SS11[31][8] = 4'h3;
    SS11[32][8] = 4'h3;
    SS11[33][8] = 4'h0;
    SS11[34][8] = 4'hD;
    SS11[35][8] = 4'hD;
    SS11[36][8] = 4'hD;
    SS11[37][8] = 4'hD;
    SS11[38][8] = 4'hD;
    SS11[39][8] = 4'hD;
    SS11[40][8] = 4'h0;
    SS11[41][8] = 4'h0;
    SS11[42][8] = 4'h0;
    SS11[43][8] = 4'h0;
    SS11[44][8] = 4'h0;
    SS11[45][8] = 4'h0;
    SS11[46][8] = 4'h0;
    SS11[47][8] = 4'h0;
    SS11[0][9] = 4'h0;
    SS11[1][9] = 4'h0;
    SS11[2][9] = 4'h0;
    SS11[3][9] = 4'h0;
    SS11[4][9] = 4'h0;
    SS11[5][9] = 4'h0;
    SS11[6][9] = 4'h0;
    SS11[7][9] = 4'h0;
    SS11[8][9] = 4'h0;
    SS11[9][9] = 4'h0;
    SS11[10][9] = 4'h0;
    SS11[11][9] = 4'h0;
    SS11[12][9] = 4'h0;
    SS11[13][9] = 4'h0;
    SS11[14][9] = 4'h0;
    SS11[15][9] = 4'h0;
    SS11[16][9] = 4'h0;
    SS11[17][9] = 4'h0;
    SS11[18][9] = 4'h0;
    SS11[19][9] = 4'h0;
    SS11[20][9] = 4'h0;
    SS11[21][9] = 4'h0;
    SS11[22][9] = 4'h0;
    SS11[23][9] = 4'h0;
    SS11[24][9] = 4'h0;
    SS11[25][9] = 4'h0;
    SS11[26][9] = 4'h0;
    SS11[27][9] = 4'h0;
    SS11[28][9] = 4'h0;
    SS11[29][9] = 4'h0;
    SS11[30][9] = 4'h3;
    SS11[31][9] = 4'h3;
    SS11[32][9] = 4'h3;
    SS11[33][9] = 4'hD;
    SS11[34][9] = 4'hD;
    SS11[35][9] = 4'hD;
    SS11[36][9] = 4'hD;
    SS11[37][9] = 4'hD;
    SS11[38][9] = 4'hD;
    SS11[39][9] = 4'hD;
    SS11[40][9] = 4'h0;
    SS11[41][9] = 4'h0;
    SS11[42][9] = 4'h0;
    SS11[43][9] = 4'h0;
    SS11[44][9] = 4'h0;
    SS11[45][9] = 4'h0;
    SS11[46][9] = 4'h0;
    SS11[47][9] = 4'h0;
    SS11[0][10] = 4'h0;
    SS11[1][10] = 4'h0;
    SS11[2][10] = 4'h0;
    SS11[3][10] = 4'h0;
    SS11[4][10] = 4'h0;
    SS11[5][10] = 4'h0;
    SS11[6][10] = 4'h0;
    SS11[7][10] = 4'h0;
    SS11[8][10] = 4'h0;
    SS11[9][10] = 4'h0;
    SS11[10][10] = 4'h0;
    SS11[11][10] = 4'h0;
    SS11[12][10] = 4'h0;
    SS11[13][10] = 4'h0;
    SS11[14][10] = 4'h0;
    SS11[15][10] = 4'h0;
    SS11[16][10] = 4'h0;
    SS11[17][10] = 4'h0;
    SS11[18][10] = 4'h0;
    SS11[19][10] = 4'h0;
    SS11[20][10] = 4'h0;
    SS11[21][10] = 4'h0;
    SS11[22][10] = 4'h0;
    SS11[23][10] = 4'h0;
    SS11[24][10] = 4'h0;
    SS11[25][10] = 4'h0;
    SS11[26][10] = 4'h0;
    SS11[27][10] = 4'h0;
    SS11[28][10] = 4'h0;
    SS11[29][10] = 4'h0;
    SS11[30][10] = 4'h3;
    SS11[31][10] = 4'h3;
    SS11[32][10] = 4'h3;
    SS11[33][10] = 4'hD;
    SS11[34][10] = 4'hD;
    SS11[35][10] = 4'hD;
    SS11[36][10] = 4'hE;
    SS11[37][10] = 4'hE;
    SS11[38][10] = 4'hD;
    SS11[39][10] = 4'h0;
    SS11[40][10] = 4'h0;
    SS11[41][10] = 4'h0;
    SS11[42][10] = 4'h0;
    SS11[43][10] = 4'h0;
    SS11[44][10] = 4'h0;
    SS11[45][10] = 4'h0;
    SS11[46][10] = 4'h0;
    SS11[47][10] = 4'h0;
    SS11[0][11] = 4'h0;
    SS11[1][11] = 4'h0;
    SS11[2][11] = 4'h0;
    SS11[3][11] = 4'h0;
    SS11[4][11] = 4'h0;
    SS11[5][11] = 4'h0;
    SS11[6][11] = 4'h0;
    SS11[7][11] = 4'h0;
    SS11[8][11] = 4'h0;
    SS11[9][11] = 4'h0;
    SS11[10][11] = 4'h0;
    SS11[11][11] = 4'h0;
    SS11[12][11] = 4'h0;
    SS11[13][11] = 4'h0;
    SS11[14][11] = 4'h0;
    SS11[15][11] = 4'h0;
    SS11[16][11] = 4'h0;
    SS11[17][11] = 4'h0;
    SS11[18][11] = 4'h0;
    SS11[19][11] = 4'h0;
    SS11[20][11] = 4'h0;
    SS11[21][11] = 4'h0;
    SS11[22][11] = 4'h0;
    SS11[23][11] = 4'h3;
    SS11[24][11] = 4'h3;
    SS11[25][11] = 4'h0;
    SS11[26][11] = 4'h0;
    SS11[27][11] = 4'h0;
    SS11[28][11] = 4'h0;
    SS11[29][11] = 4'hD;
    SS11[30][11] = 4'hD;
    SS11[31][11] = 4'hD;
    SS11[32][11] = 4'hE;
    SS11[33][11] = 4'hD;
    SS11[34][11] = 4'hD;
    SS11[35][11] = 4'hD;
    SS11[36][11] = 4'hE;
    SS11[37][11] = 4'hE;
    SS11[38][11] = 4'hE;
    SS11[39][11] = 4'h0;
    SS11[40][11] = 4'h0;
    SS11[41][11] = 4'h0;
    SS11[42][11] = 4'h0;
    SS11[43][11] = 4'h0;
    SS11[44][11] = 4'h0;
    SS11[45][11] = 4'h0;
    SS11[46][11] = 4'h0;
    SS11[47][11] = 4'h0;
    SS11[0][12] = 4'h0;
    SS11[1][12] = 4'h0;
    SS11[2][12] = 4'h0;
    SS11[3][12] = 4'hC;
    SS11[4][12] = 4'h0;
    SS11[5][12] = 4'h0;
    SS11[6][12] = 4'h0;
    SS11[7][12] = 4'h0;
    SS11[8][12] = 4'h0;
    SS11[9][12] = 4'hF;
    SS11[10][12] = 4'hD;
    SS11[11][12] = 4'hD;
    SS11[12][12] = 4'h0;
    SS11[13][12] = 4'h0;
    SS11[14][12] = 4'h0;
    SS11[15][12] = 4'h0;
    SS11[16][12] = 4'h0;
    SS11[17][12] = 4'h0;
    SS11[18][12] = 4'h0;
    SS11[19][12] = 4'h0;
    SS11[20][12] = 4'h0;
    SS11[21][12] = 4'h0;
    SS11[22][12] = 4'h3;
    SS11[23][12] = 4'h3;
    SS11[24][12] = 4'h3;
    SS11[25][12] = 4'h3;
    SS11[26][12] = 4'hD;
    SS11[27][12] = 4'h0;
    SS11[28][12] = 4'h0;
    SS11[29][12] = 4'hD;
    SS11[30][12] = 4'hD;
    SS11[31][12] = 4'hD;
    SS11[32][12] = 4'hE;
    SS11[33][12] = 4'hE;
    SS11[34][12] = 4'hE;
    SS11[35][12] = 4'hE;
    SS11[36][12] = 4'hE;
    SS11[37][12] = 4'hE;
    SS11[38][12] = 4'h0;
    SS11[39][12] = 4'h0;
    SS11[40][12] = 4'h0;
    SS11[41][12] = 4'h0;
    SS11[42][12] = 4'h0;
    SS11[43][12] = 4'h0;
    SS11[44][12] = 4'h0;
    SS11[45][12] = 4'h0;
    SS11[46][12] = 4'h0;
    SS11[47][12] = 4'h0;
    SS11[0][13] = 4'h0;
    SS11[1][13] = 4'h0;
    SS11[2][13] = 4'h0;
    SS11[3][13] = 4'hC;
    SS11[4][13] = 4'hC;
    SS11[5][13] = 4'hC;
    SS11[6][13] = 4'h0;
    SS11[7][13] = 4'h0;
    SS11[8][13] = 4'h0;
    SS11[9][13] = 4'hD;
    SS11[10][13] = 4'hD;
    SS11[11][13] = 4'hD;
    SS11[12][13] = 4'hD;
    SS11[13][13] = 4'hD;
    SS11[14][13] = 4'h0;
    SS11[15][13] = 4'h0;
    SS11[16][13] = 4'h0;
    SS11[17][13] = 4'h0;
    SS11[18][13] = 4'h0;
    SS11[19][13] = 4'h0;
    SS11[20][13] = 4'h0;
    SS11[21][13] = 4'h0;
    SS11[22][13] = 4'h3;
    SS11[23][13] = 4'h3;
    SS11[24][13] = 4'h3;
    SS11[25][13] = 4'hD;
    SS11[26][13] = 4'hD;
    SS11[27][13] = 4'hD;
    SS11[28][13] = 4'hD;
    SS11[29][13] = 4'hD;
    SS11[30][13] = 4'hD;
    SS11[31][13] = 4'hD;
    SS11[32][13] = 4'hE;
    SS11[33][13] = 4'hE;
    SS11[34][13] = 4'hE;
    SS11[35][13] = 4'hE;
    SS11[36][13] = 4'hE;
    SS11[37][13] = 4'hE;
    SS11[38][13] = 4'h0;
    SS11[39][13] = 4'h0;
    SS11[40][13] = 4'h0;
    SS11[41][13] = 4'h0;
    SS11[42][13] = 4'h0;
    SS11[43][13] = 4'h0;
    SS11[44][13] = 4'h0;
    SS11[45][13] = 4'h0;
    SS11[46][13] = 4'h0;
    SS11[47][13] = 4'h0;
    SS11[0][14] = 4'h0;
    SS11[1][14] = 4'h0;
    SS11[2][14] = 4'hC;
    SS11[3][14] = 4'hC;
    SS11[4][14] = 4'hC;
    SS11[5][14] = 4'hC;
    SS11[6][14] = 4'hC;
    SS11[7][14] = 4'hC;
    SS11[8][14] = 4'hC;
    SS11[9][14] = 4'hD;
    SS11[10][14] = 4'hD;
    SS11[11][14] = 4'hD;
    SS11[12][14] = 4'hD;
    SS11[13][14] = 4'hD;
    SS11[14][14] = 4'hD;
    SS11[15][14] = 4'hD;
    SS11[16][14] = 4'hD;
    SS11[17][14] = 4'h0;
    SS11[18][14] = 4'h0;
    SS11[19][14] = 4'h0;
    SS11[20][14] = 4'h0;
    SS11[21][14] = 4'hF;
    SS11[22][14] = 4'hD;
    SS11[23][14] = 4'hD;
    SS11[24][14] = 4'h3;
    SS11[25][14] = 4'hD;
    SS11[26][14] = 4'hD;
    SS11[27][14] = 4'hD;
    SS11[28][14] = 4'hD;
    SS11[29][14] = 4'hD;
    SS11[30][14] = 4'hD;
    SS11[31][14] = 4'hE;
    SS11[32][14] = 4'hE;
    SS11[33][14] = 4'hE;
    SS11[34][14] = 4'hE;
    SS11[35][14] = 4'hE;
    SS11[36][14] = 4'hE;
    SS11[37][14] = 4'hE;
    SS11[38][14] = 4'h0;
    SS11[39][14] = 4'h0;
    SS11[40][14] = 4'h0;
    SS11[41][14] = 4'h0;
    SS11[42][14] = 4'h0;
    SS11[43][14] = 4'h0;
    SS11[44][14] = 4'h0;
    SS11[45][14] = 4'h0;
    SS11[46][14] = 4'h0;
    SS11[47][14] = 4'h0;
    SS11[0][15] = 4'h0;
    SS11[1][15] = 4'h0;
    SS11[2][15] = 4'hC;
    SS11[3][15] = 4'hC;
    SS11[4][15] = 4'hC;
    SS11[5][15] = 4'hC;
    SS11[6][15] = 4'hC;
    SS11[7][15] = 4'hC;
    SS11[8][15] = 4'hC;
    SS11[9][15] = 4'hC;
    SS11[10][15] = 4'hC;
    SS11[11][15] = 4'hD;
    SS11[12][15] = 4'hD;
    SS11[13][15] = 4'hD;
    SS11[14][15] = 4'hD;
    SS11[15][15] = 4'hD;
    SS11[16][15] = 4'hD;
    SS11[17][15] = 4'hD;
    SS11[18][15] = 4'hC;
    SS11[19][15] = 4'h0;
    SS11[20][15] = 4'h0;
    SS11[21][15] = 4'hD;
    SS11[22][15] = 4'hD;
    SS11[23][15] = 4'hD;
    SS11[24][15] = 4'hD;
    SS11[25][15] = 4'hD;
    SS11[26][15] = 4'hD;
    SS11[27][15] = 4'hD;
    SS11[28][15] = 4'hD;
    SS11[29][15] = 4'hD;
    SS11[30][15] = 4'hD;
    SS11[31][15] = 4'hE;
    SS11[32][15] = 4'hE;
    SS11[33][15] = 4'hE;
    SS11[34][15] = 4'hE;
    SS11[35][15] = 4'hE;
    SS11[36][15] = 4'hE;
    SS11[37][15] = 4'h0;
    SS11[38][15] = 4'h0;
    SS11[39][15] = 4'h0;
    SS11[40][15] = 4'h0;
    SS11[41][15] = 4'h0;
    SS11[42][15] = 4'h0;
    SS11[43][15] = 4'h0;
    SS11[44][15] = 4'h0;
    SS11[45][15] = 4'h0;
    SS11[46][15] = 4'h0;
    SS11[47][15] = 4'h0;
    SS11[0][16] = 4'h0;
    SS11[1][16] = 4'hC;
    SS11[2][16] = 4'hC;
    SS11[3][16] = 4'hC;
    SS11[4][16] = 4'hC;
    SS11[5][16] = 4'hC;
    SS11[6][16] = 4'hC;
    SS11[7][16] = 4'hC;
    SS11[8][16] = 4'hC;
    SS11[9][16] = 4'hC;
    SS11[10][16] = 4'hC;
    SS11[11][16] = 4'hC;
    SS11[12][16] = 4'hC;
    SS11[13][16] = 4'hC;
    SS11[14][16] = 4'hD;
    SS11[15][16] = 4'hD;
    SS11[16][16] = 4'hD;
    SS11[17][16] = 4'hC;
    SS11[18][16] = 4'hC;
    SS11[19][16] = 4'hC;
    SS11[20][16] = 4'hC;
    SS11[21][16] = 4'hD;
    SS11[22][16] = 4'hD;
    SS11[23][16] = 4'hD;
    SS11[24][16] = 4'hD;
    SS11[25][16] = 4'hD;
    SS11[26][16] = 4'hD;
    SS11[27][16] = 4'hE;
    SS11[28][16] = 4'hE;
    SS11[29][16] = 4'hD;
    SS11[30][16] = 4'hE;
    SS11[31][16] = 4'hE;
    SS11[32][16] = 4'hE;
    SS11[33][16] = 4'hE;
    SS11[34][16] = 4'hC;
    SS11[35][16] = 4'hC;
    SS11[36][16] = 4'hC;
    SS11[37][16] = 4'h0;
    SS11[38][16] = 4'h0;
    SS11[39][16] = 4'h0;
    SS11[40][16] = 4'h0;
    SS11[41][16] = 4'h0;
    SS11[42][16] = 4'h0;
    SS11[43][16] = 4'hC;
    SS11[44][16] = 4'hC;
    SS11[45][16] = 4'h0;
    SS11[46][16] = 4'h0;
    SS11[47][16] = 4'h0;
    SS11[0][17] = 4'h0;
    SS11[1][17] = 4'hC;
    SS11[2][17] = 4'hC;
    SS11[3][17] = 4'hC;
    SS11[4][17] = 4'hC;
    SS11[5][17] = 4'hC;
    SS11[6][17] = 4'hC;
    SS11[7][17] = 4'hC;
    SS11[8][17] = 4'hC;
    SS11[9][17] = 4'hC;
    SS11[10][17] = 4'hC;
    SS11[11][17] = 4'hC;
    SS11[12][17] = 4'hC;
    SS11[13][17] = 4'hC;
    SS11[14][17] = 4'hC;
    SS11[15][17] = 4'hC;
    SS11[16][17] = 4'hD;
    SS11[17][17] = 4'hC;
    SS11[18][17] = 4'hC;
    SS11[19][17] = 4'hC;
    SS11[20][17] = 4'hD;
    SS11[21][17] = 4'hD;
    SS11[22][17] = 4'hD;
    SS11[23][17] = 4'hC;
    SS11[24][17] = 4'hD;
    SS11[25][17] = 4'hD;
    SS11[26][17] = 4'hD;
    SS11[27][17] = 4'hE;
    SS11[28][17] = 4'hE;
    SS11[29][17] = 4'hE;
    SS11[30][17] = 4'hC;
    SS11[31][17] = 4'hC;
    SS11[32][17] = 4'hE;
    SS11[33][17] = 4'hC;
    SS11[34][17] = 4'hC;
    SS11[35][17] = 4'hC;
    SS11[36][17] = 4'hC;
    SS11[37][17] = 4'hC;
    SS11[38][17] = 4'hC;
    SS11[39][17] = 4'h0;
    SS11[40][17] = 4'h0;
    SS11[41][17] = 4'h0;
    SS11[42][17] = 4'h0;
    SS11[43][17] = 4'hC;
    SS11[44][17] = 4'hC;
    SS11[45][17] = 4'hC;
    SS11[46][17] = 4'hC;
    SS11[47][17] = 4'h0;
    SS11[0][18] = 4'h0;
    SS11[1][18] = 4'h0;
    SS11[2][18] = 4'h0;
    SS11[3][18] = 4'hC;
    SS11[4][18] = 4'hC;
    SS11[5][18] = 4'hC;
    SS11[6][18] = 4'hC;
    SS11[7][18] = 4'hC;
    SS11[8][18] = 4'hC;
    SS11[9][18] = 4'hC;
    SS11[10][18] = 4'hC;
    SS11[11][18] = 4'hC;
    SS11[12][18] = 4'hC;
    SS11[13][18] = 4'hC;
    SS11[14][18] = 4'hC;
    SS11[15][18] = 4'hC;
    SS11[16][18] = 4'hC;
    SS11[17][18] = 4'hC;
    SS11[18][18] = 4'hC;
    SS11[19][18] = 4'hC;
    SS11[20][18] = 4'hD;
    SS11[21][18] = 4'hD;
    SS11[22][18] = 4'hD;
    SS11[23][18] = 4'hC;
    SS11[24][18] = 4'hC;
    SS11[25][18] = 4'hC;
    SS11[26][18] = 4'hE;
    SS11[27][18] = 4'hE;
    SS11[28][18] = 4'hE;
    SS11[29][18] = 4'hC;
    SS11[30][18] = 4'hC;
    SS11[31][18] = 4'hC;
    SS11[32][18] = 4'hC;
    SS11[33][18] = 4'hC;
    SS11[34][18] = 4'hC;
    SS11[35][18] = 4'hC;
    SS11[36][18] = 4'hC;
    SS11[37][18] = 4'hC;
    SS11[38][18] = 4'hC;
    SS11[39][18] = 4'hC;
    SS11[40][18] = 4'hC;
    SS11[41][18] = 4'hC;
    SS11[42][18] = 4'hC;
    SS11[43][18] = 4'hC;
    SS11[44][18] = 4'hC;
    SS11[45][18] = 4'hC;
    SS11[46][18] = 4'hC;
    SS11[47][18] = 4'hC;
    SS11[0][19] = 4'h0;
    SS11[1][19] = 4'h0;
    SS11[2][19] = 4'h0;
    SS11[3][19] = 4'h0;
    SS11[4][19] = 4'h0;
    SS11[5][19] = 4'hC;
    SS11[6][19] = 4'hC;
    SS11[7][19] = 4'hC;
    SS11[8][19] = 4'hC;
    SS11[9][19] = 4'hC;
    SS11[10][19] = 4'hC;
    SS11[11][19] = 4'hC;
    SS11[12][19] = 4'hC;
    SS11[13][19] = 4'hC;
    SS11[14][19] = 4'hC;
    SS11[15][19] = 4'hC;
    SS11[16][19] = 4'hC;
    SS11[17][19] = 4'hC;
    SS11[18][19] = 4'hC;
    SS11[19][19] = 4'hA;
    SS11[20][19] = 4'hA;
    SS11[21][19] = 4'hD;
    SS11[22][19] = 4'hD;
    SS11[23][19] = 4'hC;
    SS11[24][19] = 4'hC;
    SS11[25][19] = 4'hC;
    SS11[26][19] = 4'hC;
    SS11[27][19] = 4'hC;
    SS11[28][19] = 4'hC;
    SS11[29][19] = 4'hC;
    SS11[30][19] = 4'hC;
    SS11[31][19] = 4'hC;
    SS11[32][19] = 4'hC;
    SS11[33][19] = 4'hC;
    SS11[34][19] = 4'hC;
    SS11[35][19] = 4'hC;
    SS11[36][19] = 4'hC;
    SS11[37][19] = 4'hC;
    SS11[38][19] = 4'hC;
    SS11[39][19] = 4'hC;
    SS11[40][19] = 4'hC;
    SS11[41][19] = 4'hC;
    SS11[42][19] = 4'hC;
    SS11[43][19] = 4'hC;
    SS11[44][19] = 4'hC;
    SS11[45][19] = 4'hC;
    SS11[46][19] = 4'hC;
    SS11[47][19] = 4'hC;
    SS11[0][20] = 4'h0;
    SS11[1][20] = 4'h0;
    SS11[2][20] = 4'h0;
    SS11[3][20] = 4'h0;
    SS11[4][20] = 4'h0;
    SS11[5][20] = 4'h0;
    SS11[6][20] = 4'hD;
    SS11[7][20] = 4'hD;
    SS11[8][20] = 4'hC;
    SS11[9][20] = 4'hC;
    SS11[10][20] = 4'hC;
    SS11[11][20] = 4'hC;
    SS11[12][20] = 4'hC;
    SS11[13][20] = 4'hC;
    SS11[14][20] = 4'hC;
    SS11[15][20] = 4'hC;
    SS11[16][20] = 4'hC;
    SS11[17][20] = 4'hC;
    SS11[18][20] = 4'hC;
    SS11[19][20] = 4'hA;
    SS11[20][20] = 4'hA;
    SS11[21][20] = 4'hA;
    SS11[22][20] = 4'hD;
    SS11[23][20] = 4'hC;
    SS11[24][20] = 4'hC;
    SS11[25][20] = 4'hC;
    SS11[26][20] = 4'hC;
    SS11[27][20] = 4'hC;
    SS11[28][20] = 4'hC;
    SS11[29][20] = 4'hC;
    SS11[30][20] = 4'hC;
    SS11[31][20] = 4'hC;
    SS11[32][20] = 4'hC;
    SS11[33][20] = 4'hC;
    SS11[34][20] = 4'hC;
    SS11[35][20] = 4'hC;
    SS11[36][20] = 4'hC;
    SS11[37][20] = 4'hC;
    SS11[38][20] = 4'hD;
    SS11[39][20] = 4'hC;
    SS11[40][20] = 4'hC;
    SS11[41][20] = 4'hC;
    SS11[42][20] = 4'hC;
    SS11[43][20] = 4'hC;
    SS11[44][20] = 4'hC;
    SS11[45][20] = 4'hD;
    SS11[46][20] = 4'hD;
    SS11[47][20] = 4'hC;
    SS11[0][21] = 4'h0;
    SS11[1][21] = 4'h0;
    SS11[2][21] = 4'h0;
    SS11[3][21] = 4'h0;
    SS11[4][21] = 4'h0;
    SS11[5][21] = 4'h0;
    SS11[6][21] = 4'hD;
    SS11[7][21] = 4'hD;
    SS11[8][21] = 4'hD;
    SS11[9][21] = 4'hD;
    SS11[10][21] = 4'hC;
    SS11[11][21] = 4'hC;
    SS11[12][21] = 4'hC;
    SS11[13][21] = 4'hC;
    SS11[14][21] = 4'hC;
    SS11[15][21] = 4'hC;
    SS11[16][21] = 4'hC;
    SS11[17][21] = 4'hC;
    SS11[18][21] = 4'hC;
    SS11[19][21] = 4'hA;
    SS11[20][21] = 4'hA;
    SS11[21][21] = 4'hA;
    SS11[22][21] = 4'hD;
    SS11[23][21] = 4'hD;
    SS11[24][21] = 4'hD;
    SS11[25][21] = 4'hC;
    SS11[26][21] = 4'hC;
    SS11[27][21] = 4'hC;
    SS11[28][21] = 4'hC;
    SS11[29][21] = 4'hC;
    SS11[30][21] = 4'hC;
    SS11[31][21] = 4'hC;
    SS11[32][21] = 4'hC;
    SS11[33][21] = 4'hC;
    SS11[34][21] = 4'hC;
    SS11[35][21] = 4'hC;
    SS11[36][21] = 4'hC;
    SS11[37][21] = 4'hC;
    SS11[38][21] = 4'hD;
    SS11[39][21] = 4'hD;
    SS11[40][21] = 4'hD;
    SS11[41][21] = 4'hC;
    SS11[42][21] = 4'hC;
    SS11[43][21] = 4'hC;
    SS11[44][21] = 4'hD;
    SS11[45][21] = 4'hD;
    SS11[46][21] = 4'hD;
    SS11[47][21] = 4'h0;
    SS11[0][22] = 4'h0;
    SS11[1][22] = 4'h0;
    SS11[2][22] = 4'h0;
    SS11[3][22] = 4'h0;
    SS11[4][22] = 4'h0;
    SS11[5][22] = 4'hD;
    SS11[6][22] = 4'hD;
    SS11[7][22] = 4'hD;
    SS11[8][22] = 4'hD;
    SS11[9][22] = 4'hD;
    SS11[10][22] = 4'hD;
    SS11[11][22] = 4'hD;
    SS11[12][22] = 4'hD;
    SS11[13][22] = 4'hC;
    SS11[14][22] = 4'hC;
    SS11[15][22] = 4'hC;
    SS11[16][22] = 4'hC;
    SS11[17][22] = 4'hC;
    SS11[18][22] = 4'hA;
    SS11[19][22] = 4'hA;
    SS11[20][22] = 4'hA;
    SS11[21][22] = 4'hD;
    SS11[22][22] = 4'hD;
    SS11[23][22] = 4'hD;
    SS11[24][22] = 4'hD;
    SS11[25][22] = 4'hC;
    SS11[26][22] = 4'hC;
    SS11[27][22] = 4'hC;
    SS11[28][22] = 4'hC;
    SS11[29][22] = 4'hC;
    SS11[30][22] = 4'hC;
    SS11[31][22] = 4'hC;
    SS11[32][22] = 4'hC;
    SS11[33][22] = 4'hC;
    SS11[34][22] = 4'hD;
    SS11[35][22] = 4'hD;
    SS11[36][22] = 4'hC;
    SS11[37][22] = 4'hD;
    SS11[38][22] = 4'hD;
    SS11[39][22] = 4'hD;
    SS11[40][22] = 4'hD;
    SS11[41][22] = 4'hE;
    SS11[42][22] = 4'hE;
    SS11[43][22] = 4'hE;
    SS11[44][22] = 4'hD;
    SS11[45][22] = 4'hD;
    SS11[46][22] = 4'hD;
    SS11[47][22] = 4'h0;
    SS11[0][23] = 4'h0;
    SS11[1][23] = 4'h0;
    SS11[2][23] = 4'h0;
    SS11[3][23] = 4'h0;
    SS11[4][23] = 4'h0;
    SS11[5][23] = 4'h0;
    SS11[6][23] = 4'h0;
    SS11[7][23] = 4'hD;
    SS11[8][23] = 4'hD;
    SS11[9][23] = 4'hD;
    SS11[10][23] = 4'hD;
    SS11[11][23] = 4'hD;
    SS11[12][23] = 4'hD;
    SS11[13][23] = 4'hD;
    SS11[14][23] = 4'hD;
    SS11[15][23] = 4'hC;
    SS11[16][23] = 4'hC;
    SS11[17][23] = 4'hC;
    SS11[18][23] = 4'hA;
    SS11[19][23] = 4'hA;
    SS11[20][23] = 4'hA;
    SS11[21][23] = 4'hD;
    SS11[22][23] = 4'hD;
    SS11[23][23] = 4'hD;
    SS11[24][23] = 4'hC;
    SS11[25][23] = 4'hC;
    SS11[26][23] = 4'hC;
    SS11[27][23] = 4'hD;
    SS11[28][23] = 4'hD;
    SS11[29][23] = 4'hD;
    SS11[30][23] = 4'hD;
    SS11[31][23] = 4'hC;
    SS11[32][23] = 4'hC;
    SS11[33][23] = 4'hC;
    SS11[34][23] = 4'hD;
    SS11[35][23] = 4'hD;
    SS11[36][23] = 4'hD;
    SS11[37][23] = 4'hE;
    SS11[38][23] = 4'hD;
    SS11[39][23] = 4'hD;
    SS11[40][23] = 4'hE;
    SS11[41][23] = 4'hE;
    SS11[42][23] = 4'hE;
    SS11[43][23] = 4'h0;
    SS11[44][23] = 4'h0;
    SS11[45][23] = 4'h0;
    SS11[46][23] = 4'hD;
    SS11[47][23] = 4'h0;
    SS11[0][24] = 4'h0;
    SS11[1][24] = 4'h0;
    SS11[2][24] = 4'h0;
    SS11[3][24] = 4'h0;
    SS11[4][24] = 4'h0;
    SS11[5][24] = 4'h0;
    SS11[6][24] = 4'h0;
    SS11[7][24] = 4'h0;
    SS11[8][24] = 4'h0;
    SS11[9][24] = 4'h0;
    SS11[10][24] = 4'hD;
    SS11[11][24] = 4'hD;
    SS11[12][24] = 4'hD;
    SS11[13][24] = 4'hD;
    SS11[14][24] = 4'hC;
    SS11[15][24] = 4'hC;
    SS11[16][24] = 4'hC;
    SS11[17][24] = 4'hA;
    SS11[18][24] = 4'hA;
    SS11[19][24] = 4'hA;
    SS11[20][24] = 4'hA;
    SS11[21][24] = 4'hD;
    SS11[22][24] = 4'hD;
    SS11[23][24] = 4'hD;
    SS11[24][24] = 4'hC;
    SS11[25][24] = 4'hC;
    SS11[26][24] = 4'hC;
    SS11[27][24] = 4'hD;
    SS11[28][24] = 4'hD;
    SS11[29][24] = 4'hD;
    SS11[30][24] = 4'hE;
    SS11[31][24] = 4'hE;
    SS11[32][24] = 4'hE;
    SS11[33][24] = 4'hD;
    SS11[34][24] = 4'hD;
    SS11[35][24] = 4'hD;
    SS11[36][24] = 4'hD;
    SS11[37][24] = 4'hE;
    SS11[38][24] = 4'hE;
    SS11[39][24] = 4'hE;
    SS11[40][24] = 4'h0;
    SS11[41][24] = 4'hE;
    SS11[42][24] = 4'hE;
    SS11[43][24] = 4'h0;
    SS11[44][24] = 4'h0;
    SS11[45][24] = 4'h0;
    SS11[46][24] = 4'h0;
    SS11[47][24] = 4'h0;
    SS11[0][25] = 4'h0;
    SS11[1][25] = 4'h0;
    SS11[2][25] = 4'h0;
    SS11[3][25] = 4'h0;
    SS11[4][25] = 4'h0;
    SS11[5][25] = 4'h0;
    SS11[6][25] = 4'h0;
    SS11[7][25] = 4'h0;
    SS11[8][25] = 4'h0;
    SS11[9][25] = 4'h0;
    SS11[10][25] = 4'h0;
    SS11[11][25] = 4'h0;
    SS11[12][25] = 4'hD;
    SS11[13][25] = 4'hD;
    SS11[14][25] = 4'hC;
    SS11[15][25] = 4'hC;
    SS11[16][25] = 4'hC;
    SS11[17][25] = 4'hD;
    SS11[18][25] = 4'hD;
    SS11[19][25] = 4'hD;
    SS11[20][25] = 4'hD;
    SS11[21][25] = 4'hD;
    SS11[22][25] = 4'hD;
    SS11[23][25] = 4'hC;
    SS11[24][25] = 4'hC;
    SS11[25][25] = 4'hC;
    SS11[26][25] = 4'hC;
    SS11[27][25] = 4'hD;
    SS11[28][25] = 4'hD;
    SS11[29][25] = 4'hD;
    SS11[30][25] = 4'hE;
    SS11[31][25] = 4'hE;
    SS11[32][25] = 4'hE;
    SS11[33][25] = 4'hE;
    SS11[34][25] = 4'hE;
    SS11[35][25] = 4'hD;
    SS11[36][25] = 4'hE;
    SS11[37][25] = 4'hE;
    SS11[38][25] = 4'hE;
    SS11[39][25] = 4'h0;
    SS11[40][25] = 4'h0;
    SS11[41][25] = 4'h0;
    SS11[42][25] = 4'h0;
    SS11[43][25] = 4'h0;
    SS11[44][25] = 4'h0;
    SS11[45][25] = 4'h0;
    SS11[46][25] = 4'h0;
    SS11[47][25] = 4'h0;
    SS11[0][26] = 4'h0;
    SS11[1][26] = 4'h0;
    SS11[2][26] = 4'h0;
    SS11[3][26] = 4'h0;
    SS11[4][26] = 4'h0;
    SS11[5][26] = 4'h0;
    SS11[6][26] = 4'h0;
    SS11[7][26] = 4'h0;
    SS11[8][26] = 4'h0;
    SS11[9][26] = 4'h0;
    SS11[10][26] = 4'h0;
    SS11[11][26] = 4'h0;
    SS11[12][26] = 4'h0;
    SS11[13][26] = 4'h0;
    SS11[14][26] = 4'hE;
    SS11[15][26] = 4'hC;
    SS11[16][26] = 4'hC;
    SS11[17][26] = 4'hD;
    SS11[18][26] = 4'hD;
    SS11[19][26] = 4'hD;
    SS11[20][26] = 4'hC;
    SS11[21][26] = 4'hC;
    SS11[22][26] = 4'hD;
    SS11[23][26] = 4'hC;
    SS11[24][26] = 4'hC;
    SS11[25][26] = 4'hC;
    SS11[26][26] = 4'hD;
    SS11[27][26] = 4'hD;
    SS11[28][26] = 4'hD;
    SS11[29][26] = 4'hE;
    SS11[30][26] = 4'hE;
    SS11[31][26] = 4'hE;
    SS11[32][26] = 4'hE;
    SS11[33][26] = 4'hE;
    SS11[34][26] = 4'hE;
    SS11[35][26] = 4'hE;
    SS11[36][26] = 4'h0;
    SS11[37][26] = 4'h0;
    SS11[38][26] = 4'hE;
    SS11[39][26] = 4'h0;
    SS11[40][26] = 4'h0;
    SS11[41][26] = 4'h0;
    SS11[42][26] = 4'h0;
    SS11[43][26] = 4'h0;
    SS11[44][26] = 4'h0;
    SS11[45][26] = 4'h0;
    SS11[46][26] = 4'h0;
    SS11[47][26] = 4'h0;
    SS11[0][27] = 4'h0;
    SS11[1][27] = 4'h0;
    SS11[2][27] = 4'h0;
    SS11[3][27] = 4'h0;
    SS11[4][27] = 4'h0;
    SS11[5][27] = 4'h0;
    SS11[6][27] = 4'h0;
    SS11[7][27] = 4'h0;
    SS11[8][27] = 4'h0;
    SS11[9][27] = 4'h0;
    SS11[10][27] = 4'h0;
    SS11[11][27] = 4'h0;
    SS11[12][27] = 4'h0;
    SS11[13][27] = 4'h0;
    SS11[14][27] = 4'h0;
    SS11[15][27] = 4'h0;
    SS11[16][27] = 4'hD;
    SS11[17][27] = 4'hD;
    SS11[18][27] = 4'hD;
    SS11[19][27] = 4'hC;
    SS11[20][27] = 4'hC;
    SS11[21][27] = 4'hC;
    SS11[22][27] = 4'hC;
    SS11[23][27] = 4'hC;
    SS11[24][27] = 4'hC;
    SS11[25][27] = 4'hC;
    SS11[26][27] = 4'hD;
    SS11[27][27] = 4'hD;
    SS11[28][27] = 4'hD;
    SS11[29][27] = 4'hE;
    SS11[30][27] = 4'hE;
    SS11[31][27] = 4'hE;
    SS11[32][27] = 4'hE;
    SS11[33][27] = 4'hE;
    SS11[34][27] = 4'hE;
    SS11[35][27] = 4'h0;
    SS11[36][27] = 4'h0;
    SS11[37][27] = 4'h0;
    SS11[38][27] = 4'h0;
    SS11[39][27] = 4'h0;
    SS11[40][27] = 4'h0;
    SS11[41][27] = 4'h0;
    SS11[42][27] = 4'h0;
    SS11[43][27] = 4'h0;
    SS11[44][27] = 4'h0;
    SS11[45][27] = 4'h0;
    SS11[46][27] = 4'h0;
    SS11[47][27] = 4'h0;
    SS11[0][28] = 4'h0;
    SS11[1][28] = 4'h0;
    SS11[2][28] = 4'h0;
    SS11[3][28] = 4'h0;
    SS11[4][28] = 4'h0;
    SS11[5][28] = 4'h0;
    SS11[6][28] = 4'h0;
    SS11[7][28] = 4'h0;
    SS11[8][28] = 4'h0;
    SS11[9][28] = 4'h0;
    SS11[10][28] = 4'h0;
    SS11[11][28] = 4'h0;
    SS11[12][28] = 4'h0;
    SS11[13][28] = 4'h0;
    SS11[14][28] = 4'h0;
    SS11[15][28] = 4'h0;
    SS11[16][28] = 4'hD;
    SS11[17][28] = 4'hD;
    SS11[18][28] = 4'hD;
    SS11[19][28] = 4'hC;
    SS11[20][28] = 4'hC;
    SS11[21][28] = 4'hC;
    SS11[22][28] = 4'hC;
    SS11[23][28] = 4'hC;
    SS11[24][28] = 4'hC;
    SS11[25][28] = 4'hC;
    SS11[26][28] = 4'hC;
    SS11[27][28] = 4'hD;
    SS11[28][28] = 4'hD;
    SS11[29][28] = 4'hE;
    SS11[30][28] = 4'hE;
    SS11[31][28] = 4'hE;
    SS11[32][28] = 4'hE;
    SS11[33][28] = 4'hE;
    SS11[34][28] = 4'hE;
    SS11[35][28] = 4'h0;
    SS11[36][28] = 4'h0;
    SS11[37][28] = 4'h0;
    SS11[38][28] = 4'h0;
    SS11[39][28] = 4'h0;
    SS11[40][28] = 4'h0;
    SS11[41][28] = 4'h0;
    SS11[42][28] = 4'h0;
    SS11[43][28] = 4'h0;
    SS11[44][28] = 4'h0;
    SS11[45][28] = 4'h0;
    SS11[46][28] = 4'h0;
    SS11[47][28] = 4'h0;
    SS11[0][29] = 4'h0;
    SS11[1][29] = 4'h0;
    SS11[2][29] = 4'h0;
    SS11[3][29] = 4'h0;
    SS11[4][29] = 4'h0;
    SS11[5][29] = 4'h0;
    SS11[6][29] = 4'h0;
    SS11[7][29] = 4'h0;
    SS11[8][29] = 4'h0;
    SS11[9][29] = 4'h0;
    SS11[10][29] = 4'h0;
    SS11[11][29] = 4'h0;
    SS11[12][29] = 4'h0;
    SS11[13][29] = 4'h0;
    SS11[14][29] = 4'h0;
    SS11[15][29] = 4'hD;
    SS11[16][29] = 4'hD;
    SS11[17][29] = 4'hD;
    SS11[18][29] = 4'hD;
    SS11[19][29] = 4'hD;
    SS11[20][29] = 4'hD;
    SS11[21][29] = 4'hD;
    SS11[22][29] = 4'hC;
    SS11[23][29] = 4'hC;
    SS11[24][29] = 4'hC;
    SS11[25][29] = 4'hC;
    SS11[26][29] = 4'hC;
    SS11[27][29] = 4'hC;
    SS11[28][29] = 4'hC;
    SS11[29][29] = 4'hC;
    SS11[30][29] = 4'hE;
    SS11[31][29] = 4'hE;
    SS11[32][29] = 4'hE;
    SS11[33][29] = 4'hE;
    SS11[34][29] = 4'hE;
    SS11[35][29] = 4'h0;
    SS11[36][29] = 4'h0;
    SS11[37][29] = 4'h0;
    SS11[38][29] = 4'h0;
    SS11[39][29] = 4'h0;
    SS11[40][29] = 4'h0;
    SS11[41][29] = 4'h0;
    SS11[42][29] = 4'h0;
    SS11[43][29] = 4'h0;
    SS11[44][29] = 4'h0;
    SS11[45][29] = 4'h0;
    SS11[46][29] = 4'h0;
    SS11[47][29] = 4'h0;
    SS11[0][30] = 4'h0;
    SS11[1][30] = 4'h0;
    SS11[2][30] = 4'h0;
    SS11[3][30] = 4'h0;
    SS11[4][30] = 4'h0;
    SS11[5][30] = 4'h0;
    SS11[6][30] = 4'h0;
    SS11[7][30] = 4'h0;
    SS11[8][30] = 4'h0;
    SS11[9][30] = 4'h0;
    SS11[10][30] = 4'h0;
    SS11[11][30] = 4'h0;
    SS11[12][30] = 4'h0;
    SS11[13][30] = 4'h0;
    SS11[14][30] = 4'h0;
    SS11[15][30] = 4'h3;
    SS11[16][30] = 4'hD;
    SS11[17][30] = 4'hD;
    SS11[18][30] = 4'hD;
    SS11[19][30] = 4'hD;
    SS11[20][30] = 4'hD;
    SS11[21][30] = 4'hE;
    SS11[22][30] = 4'hE;
    SS11[23][30] = 4'hE;
    SS11[24][30] = 4'hC;
    SS11[25][30] = 4'hC;
    SS11[26][30] = 4'hC;
    SS11[27][30] = 4'hC;
    SS11[28][30] = 4'hC;
    SS11[29][30] = 4'hC;
    SS11[30][30] = 4'hC;
    SS11[31][30] = 4'hD;
    SS11[32][30] = 4'hE;
    SS11[33][30] = 4'hE;
    SS11[34][30] = 4'h0;
    SS11[35][30] = 4'h0;
    SS11[36][30] = 4'h0;
    SS11[37][30] = 4'h0;
    SS11[38][30] = 4'h0;
    SS11[39][30] = 4'h0;
    SS11[40][30] = 4'h0;
    SS11[41][30] = 4'h0;
    SS11[42][30] = 4'h0;
    SS11[43][30] = 4'h0;
    SS11[44][30] = 4'h0;
    SS11[45][30] = 4'h0;
    SS11[46][30] = 4'h0;
    SS11[47][30] = 4'h0;
    SS11[0][31] = 4'h0;
    SS11[1][31] = 4'h0;
    SS11[2][31] = 4'h0;
    SS11[3][31] = 4'h0;
    SS11[4][31] = 4'h0;
    SS11[5][31] = 4'h0;
    SS11[6][31] = 4'h0;
    SS11[7][31] = 4'h0;
    SS11[8][31] = 4'h0;
    SS11[9][31] = 4'h0;
    SS11[10][31] = 4'h0;
    SS11[11][31] = 4'h0;
    SS11[12][31] = 4'h0;
    SS11[13][31] = 4'h0;
    SS11[14][31] = 4'h3;
    SS11[15][31] = 4'h3;
    SS11[16][31] = 4'h3;
    SS11[17][31] = 4'h3;
    SS11[18][31] = 4'hD;
    SS11[19][31] = 4'hD;
    SS11[20][31] = 4'hD;
    SS11[21][31] = 4'hE;
    SS11[22][31] = 4'hE;
    SS11[23][31] = 4'hE;
    SS11[24][31] = 4'hC;
    SS11[25][31] = 4'hC;
    SS11[26][31] = 4'hC;
    SS11[27][31] = 4'hC;
    SS11[28][31] = 4'hC;
    SS11[29][31] = 4'hC;
    SS11[30][31] = 4'hC;
    SS11[31][31] = 4'hD;
    SS11[32][31] = 4'hD;
    SS11[33][31] = 4'hD;
    SS11[34][31] = 4'h0;
    SS11[35][31] = 4'h0;
    SS11[36][31] = 4'h0;
    SS11[37][31] = 4'h0;
    SS11[38][31] = 4'h0;
    SS11[39][31] = 4'h0;
    SS11[40][31] = 4'h0;
    SS11[41][31] = 4'h0;
    SS11[42][31] = 4'h0;
    SS11[43][31] = 4'h0;
    SS11[44][31] = 4'h0;
    SS11[45][31] = 4'h0;
    SS11[46][31] = 4'h0;
    SS11[47][31] = 4'h0;
    SS11[0][32] = 4'h0;
    SS11[1][32] = 4'h0;
    SS11[2][32] = 4'h0;
    SS11[3][32] = 4'h0;
    SS11[4][32] = 4'h0;
    SS11[5][32] = 4'h0;
    SS11[6][32] = 4'h0;
    SS11[7][32] = 4'h0;
    SS11[8][32] = 4'h0;
    SS11[9][32] = 4'h0;
    SS11[10][32] = 4'h0;
    SS11[11][32] = 4'h0;
    SS11[12][32] = 4'h0;
    SS11[13][32] = 4'h0;
    SS11[14][32] = 4'h3;
    SS11[15][32] = 4'h3;
    SS11[16][32] = 4'h3;
    SS11[17][32] = 4'hD;
    SS11[18][32] = 4'hD;
    SS11[19][32] = 4'hD;
    SS11[20][32] = 4'hD;
    SS11[21][32] = 4'hE;
    SS11[22][32] = 4'hE;
    SS11[23][32] = 4'hE;
    SS11[24][32] = 4'hC;
    SS11[25][32] = 4'hC;
    SS11[26][32] = 4'hC;
    SS11[27][32] = 4'hC;
    SS11[28][32] = 4'hC;
    SS11[29][32] = 4'hC;
    SS11[30][32] = 4'hD;
    SS11[31][32] = 4'hD;
    SS11[32][32] = 4'hD;
    SS11[33][32] = 4'hE;
    SS11[34][32] = 4'hE;
    SS11[35][32] = 4'hE;
    SS11[36][32] = 4'hE;
    SS11[37][32] = 4'h0;
    SS11[38][32] = 4'h0;
    SS11[39][32] = 4'h0;
    SS11[40][32] = 4'h0;
    SS11[41][32] = 4'h0;
    SS11[42][32] = 4'h0;
    SS11[43][32] = 4'h0;
    SS11[44][32] = 4'h0;
    SS11[45][32] = 4'h0;
    SS11[46][32] = 4'h0;
    SS11[47][32] = 4'h0;
    SS11[0][33] = 4'h0;
    SS11[1][33] = 4'h0;
    SS11[2][33] = 4'h0;
    SS11[3][33] = 4'h0;
    SS11[4][33] = 4'h0;
    SS11[5][33] = 4'h0;
    SS11[6][33] = 4'h0;
    SS11[7][33] = 4'h0;
    SS11[8][33] = 4'h0;
    SS11[9][33] = 4'h0;
    SS11[10][33] = 4'h0;
    SS11[11][33] = 4'h0;
    SS11[12][33] = 4'h0;
    SS11[13][33] = 4'h0;
    SS11[14][33] = 4'h0;
    SS11[15][33] = 4'h0;
    SS11[16][33] = 4'h3;
    SS11[17][33] = 4'hD;
    SS11[18][33] = 4'hD;
    SS11[19][33] = 4'hD;
    SS11[20][33] = 4'hD;
    SS11[21][33] = 4'hD;
    SS11[22][33] = 4'hD;
    SS11[23][33] = 4'hE;
    SS11[24][33] = 4'hC;
    SS11[25][33] = 4'hC;
    SS11[26][33] = 4'hC;
    SS11[27][33] = 4'hC;
    SS11[28][33] = 4'hC;
    SS11[29][33] = 4'hC;
    SS11[30][33] = 4'hC;
    SS11[31][33] = 4'hD;
    SS11[32][33] = 4'hD;
    SS11[33][33] = 4'hE;
    SS11[34][33] = 4'hE;
    SS11[35][33] = 4'hE;
    SS11[36][33] = 4'h0;
    SS11[37][33] = 4'h0;
    SS11[38][33] = 4'h0;
    SS11[39][33] = 4'h0;
    SS11[40][33] = 4'h0;
    SS11[41][33] = 4'h0;
    SS11[42][33] = 4'h0;
    SS11[43][33] = 4'h0;
    SS11[44][33] = 4'h0;
    SS11[45][33] = 4'h0;
    SS11[46][33] = 4'h0;
    SS11[47][33] = 4'h0;
    SS11[0][34] = 4'h0;
    SS11[1][34] = 4'h0;
    SS11[2][34] = 4'h0;
    SS11[3][34] = 4'h0;
    SS11[4][34] = 4'h0;
    SS11[5][34] = 4'h0;
    SS11[6][34] = 4'h0;
    SS11[7][34] = 4'h0;
    SS11[8][34] = 4'h0;
    SS11[9][34] = 4'h0;
    SS11[10][34] = 4'h0;
    SS11[11][34] = 4'h0;
    SS11[12][34] = 4'h0;
    SS11[13][34] = 4'h0;
    SS11[14][34] = 4'h0;
    SS11[15][34] = 4'h0;
    SS11[16][34] = 4'h0;
    SS11[17][34] = 4'h0;
    SS11[18][34] = 4'hD;
    SS11[19][34] = 4'hD;
    SS11[20][34] = 4'hD;
    SS11[21][34] = 4'hD;
    SS11[22][34] = 4'hD;
    SS11[23][34] = 4'hE;
    SS11[24][34] = 4'hE;
    SS11[25][34] = 4'hE;
    SS11[26][34] = 4'hC;
    SS11[27][34] = 4'hC;
    SS11[28][34] = 4'hC;
    SS11[29][34] = 4'hC;
    SS11[30][34] = 4'hC;
    SS11[31][34] = 4'hC;
    SS11[32][34] = 4'hD;
    SS11[33][34] = 4'hD;
    SS11[34][34] = 4'hE;
    SS11[35][34] = 4'hE;
    SS11[36][34] = 4'h0;
    SS11[37][34] = 4'h0;
    SS11[38][34] = 4'h0;
    SS11[39][34] = 4'h0;
    SS11[40][34] = 4'h0;
    SS11[41][34] = 4'h0;
    SS11[42][34] = 4'h0;
    SS11[43][34] = 4'h0;
    SS11[44][34] = 4'h0;
    SS11[45][34] = 4'h0;
    SS11[46][34] = 4'h0;
    SS11[47][34] = 4'h0;
    SS11[0][35] = 4'h0;
    SS11[1][35] = 4'h0;
    SS11[2][35] = 4'h0;
    SS11[3][35] = 4'h0;
    SS11[4][35] = 4'h0;
    SS11[5][35] = 4'h0;
    SS11[6][35] = 4'h0;
    SS11[7][35] = 4'h0;
    SS11[8][35] = 4'h0;
    SS11[9][35] = 4'h0;
    SS11[10][35] = 4'h0;
    SS11[11][35] = 4'h0;
    SS11[12][35] = 4'h0;
    SS11[13][35] = 4'h0;
    SS11[14][35] = 4'h0;
    SS11[15][35] = 4'h0;
    SS11[16][35] = 4'h0;
    SS11[17][35] = 4'h0;
    SS11[18][35] = 4'h0;
    SS11[19][35] = 4'hD;
    SS11[20][35] = 4'hD;
    SS11[21][35] = 4'hD;
    SS11[22][35] = 4'hE;
    SS11[23][35] = 4'hE;
    SS11[24][35] = 4'hE;
    SS11[25][35] = 4'hE;
    SS11[26][35] = 4'hC;
    SS11[27][35] = 4'hC;
    SS11[28][35] = 4'hC;
    SS11[29][35] = 4'hC;
    SS11[30][35] = 4'hC;
    SS11[31][35] = 4'hC;
    SS11[32][35] = 4'hD;
    SS11[33][35] = 4'hD;
    SS11[34][35] = 4'hD;
    SS11[35][35] = 4'hE;
    SS11[36][35] = 4'h0;
    SS11[37][35] = 4'h0;
    SS11[38][35] = 4'h0;
    SS11[39][35] = 4'h0;
    SS11[40][35] = 4'h0;
    SS11[41][35] = 4'h0;
    SS11[42][35] = 4'h0;
    SS11[43][35] = 4'h0;
    SS11[44][35] = 4'h0;
    SS11[45][35] = 4'h0;
    SS11[46][35] = 4'h0;
    SS11[47][35] = 4'h0;
    SS11[0][36] = 4'h0;
    SS11[1][36] = 4'h0;
    SS11[2][36] = 4'h0;
    SS11[3][36] = 4'h0;
    SS11[4][36] = 4'h0;
    SS11[5][36] = 4'h0;
    SS11[6][36] = 4'h0;
    SS11[7][36] = 4'h0;
    SS11[8][36] = 4'h0;
    SS11[9][36] = 4'h0;
    SS11[10][36] = 4'h0;
    SS11[11][36] = 4'h0;
    SS11[12][36] = 4'h0;
    SS11[13][36] = 4'h0;
    SS11[14][36] = 4'h0;
    SS11[15][36] = 4'h0;
    SS11[16][36] = 4'h0;
    SS11[17][36] = 4'h0;
    SS11[18][36] = 4'h0;
    SS11[19][36] = 4'hD;
    SS11[20][36] = 4'hD;
    SS11[21][36] = 4'hD;
    SS11[22][36] = 4'hE;
    SS11[23][36] = 4'hE;
    SS11[24][36] = 4'hE;
    SS11[25][36] = 4'hC;
    SS11[26][36] = 4'hC;
    SS11[27][36] = 4'hC;
    SS11[28][36] = 4'hC;
    SS11[29][36] = 4'hC;
    SS11[30][36] = 4'hC;
    SS11[31][36] = 4'hC;
    SS11[32][36] = 4'hD;
    SS11[33][36] = 4'hD;
    SS11[34][36] = 4'hD;
    SS11[35][36] = 4'hE;
    SS11[36][36] = 4'hE;
    SS11[37][36] = 4'hE;
    SS11[38][36] = 4'h0;
    SS11[39][36] = 4'h0;
    SS11[40][36] = 4'h0;
    SS11[41][36] = 4'h0;
    SS11[42][36] = 4'h0;
    SS11[43][36] = 4'h0;
    SS11[44][36] = 4'h0;
    SS11[45][36] = 4'h0;
    SS11[46][36] = 4'h0;
    SS11[47][36] = 4'h0;
    SS11[0][37] = 4'h0;
    SS11[1][37] = 4'h0;
    SS11[2][37] = 4'h0;
    SS11[3][37] = 4'h0;
    SS11[4][37] = 4'h0;
    SS11[5][37] = 4'h0;
    SS11[6][37] = 4'h0;
    SS11[7][37] = 4'h0;
    SS11[8][37] = 4'h0;
    SS11[9][37] = 4'h0;
    SS11[10][37] = 4'h0;
    SS11[11][37] = 4'h0;
    SS11[12][37] = 4'h0;
    SS11[13][37] = 4'h0;
    SS11[14][37] = 4'h0;
    SS11[15][37] = 4'h0;
    SS11[16][37] = 4'h0;
    SS11[17][37] = 4'h0;
    SS11[18][37] = 4'hD;
    SS11[19][37] = 4'hD;
    SS11[20][37] = 4'hD;
    SS11[21][37] = 4'hD;
    SS11[22][37] = 4'hE;
    SS11[23][37] = 4'hE;
    SS11[24][37] = 4'hE;
    SS11[25][37] = 4'hE;
    SS11[26][37] = 4'hC;
    SS11[27][37] = 4'hC;
    SS11[28][37] = 4'hC;
    SS11[29][37] = 4'hC;
    SS11[30][37] = 4'hC;
    SS11[31][37] = 4'hC;
    SS11[32][37] = 4'hC;
    SS11[33][37] = 4'hD;
    SS11[34][37] = 4'hE;
    SS11[35][37] = 4'hE;
    SS11[36][37] = 4'hE;
    SS11[37][37] = 4'hE;
    SS11[38][37] = 4'h0;
    SS11[39][37] = 4'h0;
    SS11[40][37] = 4'h0;
    SS11[41][37] = 4'h0;
    SS11[42][37] = 4'h0;
    SS11[43][37] = 4'h0;
    SS11[44][37] = 4'h0;
    SS11[45][37] = 4'h0;
    SS11[46][37] = 4'h0;
    SS11[47][37] = 4'h0;
    SS11[0][38] = 4'h0;
    SS11[1][38] = 4'h0;
    SS11[2][38] = 4'h0;
    SS11[3][38] = 4'h0;
    SS11[4][38] = 4'h0;
    SS11[5][38] = 4'h0;
    SS11[6][38] = 4'h0;
    SS11[7][38] = 4'h0;
    SS11[8][38] = 4'h0;
    SS11[9][38] = 4'h0;
    SS11[10][38] = 4'h0;
    SS11[11][38] = 4'h0;
    SS11[12][38] = 4'h0;
    SS11[13][38] = 4'h0;
    SS11[14][38] = 4'h0;
    SS11[15][38] = 4'h0;
    SS11[16][38] = 4'h0;
    SS11[17][38] = 4'h0;
    SS11[18][38] = 4'h3;
    SS11[19][38] = 4'h3;
    SS11[20][38] = 4'hD;
    SS11[21][38] = 4'hE;
    SS11[22][38] = 4'hE;
    SS11[23][38] = 4'hE;
    SS11[24][38] = 4'hE;
    SS11[25][38] = 4'hE;
    SS11[26][38] = 4'hE;
    SS11[27][38] = 4'hE;
    SS11[28][38] = 4'hC;
    SS11[29][38] = 4'hC;
    SS11[30][38] = 4'hC;
    SS11[31][38] = 4'hC;
    SS11[32][38] = 4'hC;
    SS11[33][38] = 4'hC;
    SS11[34][38] = 4'hC;
    SS11[35][38] = 4'hC;
    SS11[36][38] = 4'hE;
    SS11[37][38] = 4'h0;
    SS11[38][38] = 4'h0;
    SS11[39][38] = 4'h0;
    SS11[40][38] = 4'h0;
    SS11[41][38] = 4'h0;
    SS11[42][38] = 4'h0;
    SS11[43][38] = 4'h0;
    SS11[44][38] = 4'h0;
    SS11[45][38] = 4'h0;
    SS11[46][38] = 4'h0;
    SS11[47][38] = 4'h0;
    SS11[0][39] = 4'h0;
    SS11[1][39] = 4'h0;
    SS11[2][39] = 4'h0;
    SS11[3][39] = 4'h0;
    SS11[4][39] = 4'h0;
    SS11[5][39] = 4'h0;
    SS11[6][39] = 4'h0;
    SS11[7][39] = 4'h0;
    SS11[8][39] = 4'h0;
    SS11[9][39] = 4'h0;
    SS11[10][39] = 4'h0;
    SS11[11][39] = 4'h0;
    SS11[12][39] = 4'h0;
    SS11[13][39] = 4'h0;
    SS11[14][39] = 4'h0;
    SS11[15][39] = 4'h0;
    SS11[16][39] = 4'h0;
    SS11[17][39] = 4'h0;
    SS11[18][39] = 4'h3;
    SS11[19][39] = 4'h3;
    SS11[20][39] = 4'h3;
    SS11[21][39] = 4'hD;
    SS11[22][39] = 4'hD;
    SS11[23][39] = 4'hE;
    SS11[24][39] = 4'hE;
    SS11[25][39] = 4'hE;
    SS11[26][39] = 4'hE;
    SS11[27][39] = 4'h0;
    SS11[28][39] = 4'h0;
    SS11[29][39] = 4'h0;
    SS11[30][39] = 4'hC;
    SS11[31][39] = 4'hC;
    SS11[32][39] = 4'hC;
    SS11[33][39] = 4'hC;
    SS11[34][39] = 4'hC;
    SS11[35][39] = 4'hC;
    SS11[36][39] = 4'hC;
    SS11[37][39] = 4'hD;
    SS11[38][39] = 4'h0;
    SS11[39][39] = 4'h0;
    SS11[40][39] = 4'h0;
    SS11[41][39] = 4'h0;
    SS11[42][39] = 4'h0;
    SS11[43][39] = 4'h0;
    SS11[44][39] = 4'h0;
    SS11[45][39] = 4'h0;
    SS11[46][39] = 4'h0;
    SS11[47][39] = 4'h0;
    SS11[0][40] = 4'h0;
    SS11[1][40] = 4'h0;
    SS11[2][40] = 4'h0;
    SS11[3][40] = 4'h0;
    SS11[4][40] = 4'h0;
    SS11[5][40] = 4'h0;
    SS11[6][40] = 4'h0;
    SS11[7][40] = 4'h0;
    SS11[8][40] = 4'h0;
    SS11[9][40] = 4'h0;
    SS11[10][40] = 4'h0;
    SS11[11][40] = 4'h0;
    SS11[12][40] = 4'h0;
    SS11[13][40] = 4'h0;
    SS11[14][40] = 4'h0;
    SS11[15][40] = 4'h0;
    SS11[16][40] = 4'h0;
    SS11[17][40] = 4'h3;
    SS11[18][40] = 4'h3;
    SS11[19][40] = 4'h3;
    SS11[20][40] = 4'hD;
    SS11[21][40] = 4'hD;
    SS11[22][40] = 4'hD;
    SS11[23][40] = 4'hD;
    SS11[24][40] = 4'hE;
    SS11[25][40] = 4'hE;
    SS11[26][40] = 4'hE;
    SS11[27][40] = 4'h0;
    SS11[28][40] = 4'h0;
    SS11[29][40] = 4'h0;
    SS11[30][40] = 4'h0;
    SS11[31][40] = 4'h0;
    SS11[32][40] = 4'h0;
    SS11[33][40] = 4'hC;
    SS11[34][40] = 4'hC;
    SS11[35][40] = 4'hC;
    SS11[36][40] = 4'hD;
    SS11[37][40] = 4'hD;
    SS11[38][40] = 4'hD;
    SS11[39][40] = 4'hD;
    SS11[40][40] = 4'h0;
    SS11[41][40] = 4'h0;
    SS11[42][40] = 4'h0;
    SS11[43][40] = 4'h0;
    SS11[44][40] = 4'h0;
    SS11[45][40] = 4'h0;
    SS11[46][40] = 4'h0;
    SS11[47][40] = 4'h0;
    SS11[0][41] = 4'h0;
    SS11[1][41] = 4'h0;
    SS11[2][41] = 4'h0;
    SS11[3][41] = 4'h0;
    SS11[4][41] = 4'h0;
    SS11[5][41] = 4'h0;
    SS11[6][41] = 4'h0;
    SS11[7][41] = 4'h0;
    SS11[8][41] = 4'h0;
    SS11[9][41] = 4'h0;
    SS11[10][41] = 4'h0;
    SS11[11][41] = 4'h0;
    SS11[12][41] = 4'h0;
    SS11[13][41] = 4'h0;
    SS11[14][41] = 4'h0;
    SS11[15][41] = 4'h0;
    SS11[16][41] = 4'h0;
    SS11[17][41] = 4'h0;
    SS11[18][41] = 4'h0;
    SS11[19][41] = 4'h0;
    SS11[20][41] = 4'hD;
    SS11[21][41] = 4'hD;
    SS11[22][41] = 4'hD;
    SS11[23][41] = 4'hE;
    SS11[24][41] = 4'hE;
    SS11[25][41] = 4'hE;
    SS11[26][41] = 4'h0;
    SS11[27][41] = 4'h0;
    SS11[28][41] = 4'h0;
    SS11[29][41] = 4'h0;
    SS11[30][41] = 4'h0;
    SS11[31][41] = 4'h0;
    SS11[32][41] = 4'h0;
    SS11[33][41] = 4'hC;
    SS11[34][41] = 4'hC;
    SS11[35][41] = 4'hC;
    SS11[36][41] = 4'hD;
    SS11[37][41] = 4'hD;
    SS11[38][41] = 4'hD;
    SS11[39][41] = 4'h0;
    SS11[40][41] = 4'h0;
    SS11[41][41] = 4'h0;
    SS11[42][41] = 4'h0;
    SS11[43][41] = 4'h0;
    SS11[44][41] = 4'h0;
    SS11[45][41] = 4'h0;
    SS11[46][41] = 4'h0;
    SS11[47][41] = 4'h0;
    SS11[0][42] = 4'h0;
    SS11[1][42] = 4'h0;
    SS11[2][42] = 4'h0;
    SS11[3][42] = 4'h0;
    SS11[4][42] = 4'h0;
    SS11[5][42] = 4'h0;
    SS11[6][42] = 4'h0;
    SS11[7][42] = 4'h0;
    SS11[8][42] = 4'h0;
    SS11[9][42] = 4'h0;
    SS11[10][42] = 4'h0;
    SS11[11][42] = 4'h0;
    SS11[12][42] = 4'h0;
    SS11[13][42] = 4'h0;
    SS11[14][42] = 4'h0;
    SS11[15][42] = 4'h0;
    SS11[16][42] = 4'h0;
    SS11[17][42] = 4'h0;
    SS11[18][42] = 4'h0;
    SS11[19][42] = 4'h0;
    SS11[20][42] = 4'hD;
    SS11[21][42] = 4'hD;
    SS11[22][42] = 4'hD;
    SS11[23][42] = 4'hE;
    SS11[24][42] = 4'hE;
    SS11[25][42] = 4'hE;
    SS11[26][42] = 4'h0;
    SS11[27][42] = 4'h0;
    SS11[28][42] = 4'h0;
    SS11[29][42] = 4'h0;
    SS11[30][42] = 4'h0;
    SS11[31][42] = 4'h0;
    SS11[32][42] = 4'hC;
    SS11[33][42] = 4'hC;
    SS11[34][42] = 4'hC;
    SS11[35][42] = 4'hC;
    SS11[36][42] = 4'hC;
    SS11[37][42] = 4'hC;
    SS11[38][42] = 4'hD;
    SS11[39][42] = 4'h0;
    SS11[40][42] = 4'h0;
    SS11[41][42] = 4'h0;
    SS11[42][42] = 4'h0;
    SS11[43][42] = 4'h0;
    SS11[44][42] = 4'h0;
    SS11[45][42] = 4'h0;
    SS11[46][42] = 4'h0;
    SS11[47][42] = 4'h0;
    SS11[0][43] = 4'h0;
    SS11[1][43] = 4'h0;
    SS11[2][43] = 4'h0;
    SS11[3][43] = 4'h0;
    SS11[4][43] = 4'h0;
    SS11[5][43] = 4'h0;
    SS11[6][43] = 4'h0;
    SS11[7][43] = 4'h0;
    SS11[8][43] = 4'h0;
    SS11[9][43] = 4'h0;
    SS11[10][43] = 4'h0;
    SS11[11][43] = 4'h0;
    SS11[12][43] = 4'h0;
    SS11[13][43] = 4'h0;
    SS11[14][43] = 4'h0;
    SS11[15][43] = 4'h0;
    SS11[16][43] = 4'h0;
    SS11[17][43] = 4'h0;
    SS11[18][43] = 4'h0;
    SS11[19][43] = 4'hD;
    SS11[20][43] = 4'hD;
    SS11[21][43] = 4'hD;
    SS11[22][43] = 4'hD;
    SS11[23][43] = 4'hD;
    SS11[24][43] = 4'hD;
    SS11[25][43] = 4'hE;
    SS11[26][43] = 4'h0;
    SS11[27][43] = 4'h0;
    SS11[28][43] = 4'h0;
    SS11[29][43] = 4'h0;
    SS11[30][43] = 4'h0;
    SS11[31][43] = 4'h0;
    SS11[32][43] = 4'hC;
    SS11[33][43] = 4'hC;
    SS11[34][43] = 4'hC;
    SS11[35][43] = 4'hC;
    SS11[36][43] = 4'hC;
    SS11[37][43] = 4'hC;
    SS11[38][43] = 4'hD;
    SS11[39][43] = 4'hD;
    SS11[40][43] = 4'h0;
    SS11[41][43] = 4'h0;
    SS11[42][43] = 4'h0;
    SS11[43][43] = 4'h0;
    SS11[44][43] = 4'h0;
    SS11[45][43] = 4'h0;
    SS11[46][43] = 4'h0;
    SS11[47][43] = 4'h0;
    SS11[0][44] = 4'h0;
    SS11[1][44] = 4'h0;
    SS11[2][44] = 4'h0;
    SS11[3][44] = 4'h0;
    SS11[4][44] = 4'h0;
    SS11[5][44] = 4'h0;
    SS11[6][44] = 4'h0;
    SS11[7][44] = 4'h0;
    SS11[8][44] = 4'h0;
    SS11[9][44] = 4'h0;
    SS11[10][44] = 4'h0;
    SS11[11][44] = 4'h0;
    SS11[12][44] = 4'h0;
    SS11[13][44] = 4'h0;
    SS11[14][44] = 4'h0;
    SS11[15][44] = 4'h0;
    SS11[16][44] = 4'h0;
    SS11[17][44] = 4'h0;
    SS11[18][44] = 4'h0;
    SS11[19][44] = 4'hD;
    SS11[20][44] = 4'hD;
    SS11[21][44] = 4'hD;
    SS11[22][44] = 4'hD;
    SS11[23][44] = 4'hD;
    SS11[24][44] = 4'hD;
    SS11[25][44] = 4'h0;
    SS11[26][44] = 4'h0;
    SS11[27][44] = 4'h0;
    SS11[28][44] = 4'h0;
    SS11[29][44] = 4'h0;
    SS11[30][44] = 4'h0;
    SS11[31][44] = 4'h0;
    SS11[32][44] = 4'h0;
    SS11[33][44] = 4'h0;
    SS11[34][44] = 4'h0;
    SS11[35][44] = 4'hC;
    SS11[36][44] = 4'hC;
    SS11[37][44] = 4'hC;
    SS11[38][44] = 4'hD;
    SS11[39][44] = 4'hD;
    SS11[40][44] = 4'hD;
    SS11[41][44] = 4'h0;
    SS11[42][44] = 4'h0;
    SS11[43][44] = 4'h0;
    SS11[44][44] = 4'h0;
    SS11[45][44] = 4'h0;
    SS11[46][44] = 4'h0;
    SS11[47][44] = 4'h0;
    SS11[0][45] = 4'h0;
    SS11[1][45] = 4'h0;
    SS11[2][45] = 4'h0;
    SS11[3][45] = 4'h0;
    SS11[4][45] = 4'h0;
    SS11[5][45] = 4'h0;
    SS11[6][45] = 4'h0;
    SS11[7][45] = 4'h0;
    SS11[8][45] = 4'h0;
    SS11[9][45] = 4'h0;
    SS11[10][45] = 4'h0;
    SS11[11][45] = 4'h0;
    SS11[12][45] = 4'h0;
    SS11[13][45] = 4'h0;
    SS11[14][45] = 4'h0;
    SS11[15][45] = 4'h0;
    SS11[16][45] = 4'h0;
    SS11[17][45] = 4'h0;
    SS11[18][45] = 4'h0;
    SS11[19][45] = 4'h0;
    SS11[20][45] = 4'h0;
    SS11[21][45] = 4'hE;
    SS11[22][45] = 4'hD;
    SS11[23][45] = 4'hD;
    SS11[24][45] = 4'hD;
    SS11[25][45] = 4'h0;
    SS11[26][45] = 4'h0;
    SS11[27][45] = 4'h0;
    SS11[28][45] = 4'h0;
    SS11[29][45] = 4'h0;
    SS11[30][45] = 4'h0;
    SS11[31][45] = 4'h0;
    SS11[32][45] = 4'h0;
    SS11[33][45] = 4'h0;
    SS11[34][45] = 4'h0;
    SS11[35][45] = 4'h0;
    SS11[36][45] = 4'h0;
    SS11[37][45] = 4'hC;
    SS11[38][45] = 4'hD;
    SS11[39][45] = 4'hD;
    SS11[40][45] = 4'hD;
    SS11[41][45] = 4'h0;
    SS11[42][45] = 4'h0;
    SS11[43][45] = 4'h0;
    SS11[44][45] = 4'h0;
    SS11[45][45] = 4'h0;
    SS11[46][45] = 4'h0;
    SS11[47][45] = 4'h0;
    SS11[0][46] = 4'h0;
    SS11[1][46] = 4'h0;
    SS11[2][46] = 4'h0;
    SS11[3][46] = 4'h0;
    SS11[4][46] = 4'h0;
    SS11[5][46] = 4'h0;
    SS11[6][46] = 4'h0;
    SS11[7][46] = 4'h0;
    SS11[8][46] = 4'h0;
    SS11[9][46] = 4'h0;
    SS11[10][46] = 4'h0;
    SS11[11][46] = 4'h0;
    SS11[12][46] = 4'h0;
    SS11[13][46] = 4'h0;
    SS11[14][46] = 4'h0;
    SS11[15][46] = 4'h0;
    SS11[16][46] = 4'h0;
    SS11[17][46] = 4'h0;
    SS11[18][46] = 4'h0;
    SS11[19][46] = 4'h0;
    SS11[20][46] = 4'h0;
    SS11[21][46] = 4'hD;
    SS11[22][46] = 4'hD;
    SS11[23][46] = 4'hD;
    SS11[24][46] = 4'h0;
    SS11[25][46] = 4'h0;
    SS11[26][46] = 4'h0;
    SS11[27][46] = 4'h0;
    SS11[28][46] = 4'h0;
    SS11[29][46] = 4'h0;
    SS11[30][46] = 4'h0;
    SS11[31][46] = 4'h0;
    SS11[32][46] = 4'h0;
    SS11[33][46] = 4'h0;
    SS11[34][46] = 4'h0;
    SS11[35][46] = 4'h0;
    SS11[36][46] = 4'h0;
    SS11[37][46] = 4'h0;
    SS11[38][46] = 4'h0;
    SS11[39][46] = 4'h0;
    SS11[40][46] = 4'h0;
    SS11[41][46] = 4'h0;
    SS11[42][46] = 4'h0;
    SS11[43][46] = 4'h0;
    SS11[44][46] = 4'h0;
    SS11[45][46] = 4'h0;
    SS11[46][46] = 4'h0;
    SS11[47][46] = 4'h0;
    SS11[0][47] = 4'h0;
    SS11[1][47] = 4'h0;
    SS11[2][47] = 4'h0;
    SS11[3][47] = 4'h0;
    SS11[4][47] = 4'h0;
    SS11[5][47] = 4'h0;
    SS11[6][47] = 4'h0;
    SS11[7][47] = 4'h0;
    SS11[8][47] = 4'h0;
    SS11[9][47] = 4'h0;
    SS11[10][47] = 4'h0;
    SS11[11][47] = 4'h0;
    SS11[12][47] = 4'h0;
    SS11[13][47] = 4'h0;
    SS11[14][47] = 4'h0;
    SS11[15][47] = 4'h0;
    SS11[16][47] = 4'h0;
    SS11[17][47] = 4'h0;
    SS11[18][47] = 4'h0;
    SS11[19][47] = 4'h0;
    SS11[20][47] = 4'h0;
    SS11[21][47] = 4'hD;
    SS11[22][47] = 4'hD;
    SS11[23][47] = 4'hD;
    SS11[24][47] = 4'h0;
    SS11[25][47] = 4'h0;
    SS11[26][47] = 4'h0;
    SS11[27][47] = 4'h0;
    SS11[28][47] = 4'h0;
    SS11[29][47] = 4'h0;
    SS11[30][47] = 4'h0;
    SS11[31][47] = 4'h0;
    SS11[32][47] = 4'h0;
    SS11[33][47] = 4'h0;
    SS11[34][47] = 4'h0;
    SS11[35][47] = 4'h0;
    SS11[36][47] = 4'h0;
    SS11[37][47] = 4'h0;
    SS11[38][47] = 4'h0;
    SS11[39][47] = 4'h0;
    SS11[40][47] = 4'h0;
    SS11[41][47] = 4'h0;
    SS11[42][47] = 4'h0;
    SS11[43][47] = 4'h0;
    SS11[44][47] = 4'h0;
    SS11[45][47] = 4'h0;
    SS11[46][47] = 4'h0;
    SS11[47][47] = 4'h0;
 
//SS 12
    SS12[0][0] = 4'h0;
    SS12[1][0] = 4'h0;
    SS12[2][0] = 4'h0;
    SS12[3][0] = 4'h0;
    SS12[4][0] = 4'h0;
    SS12[5][0] = 4'h0;
    SS12[6][0] = 4'h0;
    SS12[7][0] = 4'h0;
    SS12[8][0] = 4'h0;
    SS12[9][0] = 4'h0;
    SS12[10][0] = 4'h0;
    SS12[11][0] = 4'h0;
    SS12[12][0] = 4'h0;
    SS12[13][0] = 4'h0;
    SS12[14][0] = 4'h0;
    SS12[15][0] = 4'h0;
    SS12[16][0] = 4'h0;
    SS12[17][0] = 4'h0;
    SS12[18][0] = 4'h0;
    SS12[19][0] = 4'h0;
    SS12[20][0] = 4'h0;
    SS12[21][0] = 4'h0;
    SS12[22][0] = 4'h0;
    SS12[23][0] = 4'h0;
    SS12[24][0] = 4'h0;
    SS12[25][0] = 4'h0;
    SS12[26][0] = 4'h0;
    SS12[27][0] = 4'h0;
    SS12[28][0] = 4'h0;
    SS12[29][0] = 4'h0;
    SS12[30][0] = 4'h0;
    SS12[31][0] = 4'h0;
    SS12[32][0] = 4'h0;
    SS12[33][0] = 4'h0;
    SS12[34][0] = 4'h0;
    SS12[35][0] = 4'h0;
    SS12[36][0] = 4'h0;
    SS12[37][0] = 4'h0;
    SS12[38][0] = 4'h0;
    SS12[39][0] = 4'h0;
    SS12[40][0] = 4'h0;
    SS12[41][0] = 4'h0;
    SS12[42][0] = 4'h0;
    SS12[43][0] = 4'h0;
    SS12[44][0] = 4'h0;
    SS12[45][0] = 4'h0;
    SS12[46][0] = 4'h0;
    SS12[47][0] = 4'h0;
    SS12[0][1] = 4'h0;
    SS12[1][1] = 4'h0;
    SS12[2][1] = 4'h0;
    SS12[3][1] = 4'h0;
    SS12[4][1] = 4'h0;
    SS12[5][1] = 4'h0;
    SS12[6][1] = 4'h0;
    SS12[7][1] = 4'h0;
    SS12[8][1] = 4'h0;
    SS12[9][1] = 4'h0;
    SS12[10][1] = 4'h0;
    SS12[11][1] = 4'h0;
    SS12[12][1] = 4'h0;
    SS12[13][1] = 4'h0;
    SS12[14][1] = 4'h0;
    SS12[15][1] = 4'h0;
    SS12[16][1] = 4'h0;
    SS12[17][1] = 4'h0;
    SS12[18][1] = 4'h0;
    SS12[19][1] = 4'h0;
    SS12[20][1] = 4'h0;
    SS12[21][1] = 4'h0;
    SS12[22][1] = 4'h0;
    SS12[23][1] = 4'h0;
    SS12[24][1] = 4'h0;
    SS12[25][1] = 4'h0;
    SS12[26][1] = 4'h0;
    SS12[27][1] = 4'h0;
    SS12[28][1] = 4'h0;
    SS12[29][1] = 4'h0;
    SS12[30][1] = 4'h0;
    SS12[31][1] = 4'h0;
    SS12[32][1] = 4'h0;
    SS12[33][1] = 4'h0;
    SS12[34][1] = 4'h0;
    SS12[35][1] = 4'h0;
    SS12[36][1] = 4'h0;
    SS12[37][1] = 4'h0;
    SS12[38][1] = 4'h0;
    SS12[39][1] = 4'h0;
    SS12[40][1] = 4'h0;
    SS12[41][1] = 4'h0;
    SS12[42][1] = 4'h0;
    SS12[43][1] = 4'h0;
    SS12[44][1] = 4'h0;
    SS12[45][1] = 4'h0;
    SS12[46][1] = 4'h0;
    SS12[47][1] = 4'h0;
    SS12[0][2] = 4'h0;
    SS12[1][2] = 4'h0;
    SS12[2][2] = 4'h0;
    SS12[3][2] = 4'h0;
    SS12[4][2] = 4'h0;
    SS12[5][2] = 4'h0;
    SS12[6][2] = 4'h0;
    SS12[7][2] = 4'h0;
    SS12[8][2] = 4'h0;
    SS12[9][2] = 4'h0;
    SS12[10][2] = 4'h0;
    SS12[11][2] = 4'h0;
    SS12[12][2] = 4'h0;
    SS12[13][2] = 4'h0;
    SS12[14][2] = 4'h0;
    SS12[15][2] = 4'h0;
    SS12[16][2] = 4'h0;
    SS12[17][2] = 4'h0;
    SS12[18][2] = 4'h0;
    SS12[19][2] = 4'h0;
    SS12[20][2] = 4'h0;
    SS12[21][2] = 4'h0;
    SS12[22][2] = 4'h0;
    SS12[23][2] = 4'h0;
    SS12[24][2] = 4'h0;
    SS12[25][2] = 4'h0;
    SS12[26][2] = 4'h0;
    SS12[27][2] = 4'h0;
    SS12[28][2] = 4'h0;
    SS12[29][2] = 4'h0;
    SS12[30][2] = 4'h0;
    SS12[31][2] = 4'h0;
    SS12[32][2] = 4'h0;
    SS12[33][2] = 4'h0;
    SS12[34][2] = 4'h0;
    SS12[35][2] = 4'h0;
    SS12[36][2] = 4'h0;
    SS12[37][2] = 4'h0;
    SS12[38][2] = 4'h0;
    SS12[39][2] = 4'h0;
    SS12[40][2] = 4'h0;
    SS12[41][2] = 4'h0;
    SS12[42][2] = 4'h0;
    SS12[43][2] = 4'h0;
    SS12[44][2] = 4'h0;
    SS12[45][2] = 4'h0;
    SS12[46][2] = 4'h0;
    SS12[47][2] = 4'h0;
    SS12[0][3] = 4'h0;
    SS12[1][3] = 4'h0;
    SS12[2][3] = 4'h0;
    SS12[3][3] = 4'h0;
    SS12[4][3] = 4'h0;
    SS12[5][3] = 4'h0;
    SS12[6][3] = 4'h0;
    SS12[7][3] = 4'h0;
    SS12[8][3] = 4'h0;
    SS12[9][3] = 4'h0;
    SS12[10][3] = 4'h0;
    SS12[11][3] = 4'h0;
    SS12[12][3] = 4'h0;
    SS12[13][3] = 4'h0;
    SS12[14][3] = 4'h0;
    SS12[15][3] = 4'h0;
    SS12[16][3] = 4'h0;
    SS12[17][3] = 4'h0;
    SS12[18][3] = 4'h0;
    SS12[19][3] = 4'h0;
    SS12[20][3] = 4'h0;
    SS12[21][3] = 4'h0;
    SS12[22][3] = 4'h0;
    SS12[23][3] = 4'h0;
    SS12[24][3] = 4'h0;
    SS12[25][3] = 4'h0;
    SS12[26][3] = 4'h0;
    SS12[27][3] = 4'h0;
    SS12[28][3] = 4'h0;
    SS12[29][3] = 4'h0;
    SS12[30][3] = 4'h0;
    SS12[31][3] = 4'h0;
    SS12[32][3] = 4'h0;
    SS12[33][3] = 4'h0;
    SS12[34][3] = 4'h0;
    SS12[35][3] = 4'h0;
    SS12[36][3] = 4'h0;
    SS12[37][3] = 4'h0;
    SS12[38][3] = 4'h0;
    SS12[39][3] = 4'h0;
    SS12[40][3] = 4'h0;
    SS12[41][3] = 4'h0;
    SS12[42][3] = 4'h0;
    SS12[43][3] = 4'h0;
    SS12[44][3] = 4'h0;
    SS12[45][3] = 4'h0;
    SS12[46][3] = 4'h0;
    SS12[47][3] = 4'h0;
    SS12[0][4] = 4'h0;
    SS12[1][4] = 4'h0;
    SS12[2][4] = 4'h0;
    SS12[3][4] = 4'h0;
    SS12[4][4] = 4'h0;
    SS12[5][4] = 4'h0;
    SS12[6][4] = 4'h0;
    SS12[7][4] = 4'h0;
    SS12[8][4] = 4'h0;
    SS12[9][4] = 4'h0;
    SS12[10][4] = 4'h0;
    SS12[11][4] = 4'h0;
    SS12[12][4] = 4'h0;
    SS12[13][4] = 4'h0;
    SS12[14][4] = 4'h0;
    SS12[15][4] = 4'h0;
    SS12[16][4] = 4'h0;
    SS12[17][4] = 4'h0;
    SS12[18][4] = 4'h0;
    SS12[19][4] = 4'h0;
    SS12[20][4] = 4'h0;
    SS12[21][4] = 4'h0;
    SS12[22][4] = 4'h0;
    SS12[23][4] = 4'h0;
    SS12[24][4] = 4'h0;
    SS12[25][4] = 4'h0;
    SS12[26][4] = 4'h0;
    SS12[27][4] = 4'h0;
    SS12[28][4] = 4'h0;
    SS12[29][4] = 4'h0;
    SS12[30][4] = 4'h0;
    SS12[31][4] = 4'h0;
    SS12[32][4] = 4'h0;
    SS12[33][4] = 4'h0;
    SS12[34][4] = 4'h0;
    SS12[35][4] = 4'h0;
    SS12[36][4] = 4'h0;
    SS12[37][4] = 4'h0;
    SS12[38][4] = 4'h0;
    SS12[39][4] = 4'h0;
    SS12[40][4] = 4'h0;
    SS12[41][4] = 4'h0;
    SS12[42][4] = 4'h0;
    SS12[43][4] = 4'h0;
    SS12[44][4] = 4'h0;
    SS12[45][4] = 4'h0;
    SS12[46][4] = 4'h0;
    SS12[47][4] = 4'h0;
    SS12[0][5] = 4'h0;
    SS12[1][5] = 4'h0;
    SS12[2][5] = 4'h0;
    SS12[3][5] = 4'h0;
    SS12[4][5] = 4'h0;
    SS12[5][5] = 4'h0;
    SS12[6][5] = 4'h0;
    SS12[7][5] = 4'h0;
    SS12[8][5] = 4'h0;
    SS12[9][5] = 4'hC;
    SS12[10][5] = 4'h0;
    SS12[11][5] = 4'h0;
    SS12[12][5] = 4'h0;
    SS12[13][5] = 4'h0;
    SS12[14][5] = 4'h0;
    SS12[15][5] = 4'h0;
    SS12[16][5] = 4'h0;
    SS12[17][5] = 4'h0;
    SS12[18][5] = 4'h0;
    SS12[19][5] = 4'h0;
    SS12[20][5] = 4'h0;
    SS12[21][5] = 4'h0;
    SS12[22][5] = 4'h0;
    SS12[23][5] = 4'h0;
    SS12[24][5] = 4'h0;
    SS12[25][5] = 4'h0;
    SS12[26][5] = 4'h0;
    SS12[27][5] = 4'h0;
    SS12[28][5] = 4'h0;
    SS12[29][5] = 4'h0;
    SS12[30][5] = 4'h0;
    SS12[31][5] = 4'h0;
    SS12[32][5] = 4'h0;
    SS12[33][5] = 4'h0;
    SS12[34][5] = 4'h0;
    SS12[35][5] = 4'h0;
    SS12[36][5] = 4'h0;
    SS12[37][5] = 4'h0;
    SS12[38][5] = 4'h0;
    SS12[39][5] = 4'h0;
    SS12[40][5] = 4'h0;
    SS12[41][5] = 4'h0;
    SS12[42][5] = 4'h0;
    SS12[43][5] = 4'h0;
    SS12[44][5] = 4'h0;
    SS12[45][5] = 4'h0;
    SS12[46][5] = 4'h0;
    SS12[47][5] = 4'h0;
    SS12[0][6] = 4'h0;
    SS12[1][6] = 4'h0;
    SS12[2][6] = 4'h0;
    SS12[3][6] = 4'h0;
    SS12[4][6] = 4'h0;
    SS12[5][6] = 4'h0;
    SS12[6][6] = 4'h0;
    SS12[7][6] = 4'h0;
    SS12[8][6] = 4'hC;
    SS12[9][6] = 4'hC;
    SS12[10][6] = 4'hC;
    SS12[11][6] = 4'h0;
    SS12[12][6] = 4'h0;
    SS12[13][6] = 4'h0;
    SS12[14][6] = 4'h0;
    SS12[15][6] = 4'h0;
    SS12[16][6] = 4'h0;
    SS12[17][6] = 4'h0;
    SS12[18][6] = 4'h0;
    SS12[19][6] = 4'h0;
    SS12[20][6] = 4'h0;
    SS12[21][6] = 4'h0;
    SS12[22][6] = 4'h0;
    SS12[23][6] = 4'h0;
    SS12[24][6] = 4'h0;
    SS12[25][6] = 4'h0;
    SS12[26][6] = 4'h0;
    SS12[27][6] = 4'h0;
    SS12[28][6] = 4'h0;
    SS12[29][6] = 4'h0;
    SS12[30][6] = 4'h0;
    SS12[31][6] = 4'h0;
    SS12[32][6] = 4'h0;
    SS12[33][6] = 4'h0;
    SS12[34][6] = 4'h0;
    SS12[35][6] = 4'h0;
    SS12[36][6] = 4'h0;
    SS12[37][6] = 4'h0;
    SS12[38][6] = 4'h0;
    SS12[39][6] = 4'h0;
    SS12[40][6] = 4'h0;
    SS12[41][6] = 4'h0;
    SS12[42][6] = 4'h0;
    SS12[43][6] = 4'h0;
    SS12[44][6] = 4'h0;
    SS12[45][6] = 4'h0;
    SS12[46][6] = 4'h0;
    SS12[47][6] = 4'h0;
    SS12[0][7] = 4'h0;
    SS12[1][7] = 4'h0;
    SS12[2][7] = 4'h0;
    SS12[3][7] = 4'h0;
    SS12[4][7] = 4'h0;
    SS12[5][7] = 4'h0;
    SS12[6][7] = 4'h0;
    SS12[7][7] = 4'hC;
    SS12[8][7] = 4'hC;
    SS12[9][7] = 4'hC;
    SS12[10][7] = 4'hC;
    SS12[11][7] = 4'hC;
    SS12[12][7] = 4'h0;
    SS12[13][7] = 4'h0;
    SS12[14][7] = 4'h0;
    SS12[15][7] = 4'hD;
    SS12[16][7] = 4'h0;
    SS12[17][7] = 4'h0;
    SS12[18][7] = 4'h0;
    SS12[19][7] = 4'h0;
    SS12[20][7] = 4'h0;
    SS12[21][7] = 4'h0;
    SS12[22][7] = 4'h0;
    SS12[23][7] = 4'h0;
    SS12[24][7] = 4'h0;
    SS12[25][7] = 4'h0;
    SS12[26][7] = 4'h0;
    SS12[27][7] = 4'h0;
    SS12[28][7] = 4'h0;
    SS12[29][7] = 4'h0;
    SS12[30][7] = 4'h0;
    SS12[31][7] = 4'h0;
    SS12[32][7] = 4'h0;
    SS12[33][7] = 4'h0;
    SS12[34][7] = 4'h0;
    SS12[35][7] = 4'h0;
    SS12[36][7] = 4'h0;
    SS12[37][7] = 4'h0;
    SS12[38][7] = 4'h0;
    SS12[39][7] = 4'h0;
    SS12[40][7] = 4'h0;
    SS12[41][7] = 4'h0;
    SS12[42][7] = 4'h0;
    SS12[43][7] = 4'h0;
    SS12[44][7] = 4'h0;
    SS12[45][7] = 4'h0;
    SS12[46][7] = 4'h0;
    SS12[47][7] = 4'h0;
    SS12[0][8] = 4'h0;
    SS12[1][8] = 4'h0;
    SS12[2][8] = 4'h0;
    SS12[3][8] = 4'h0;
    SS12[4][8] = 4'h0;
    SS12[5][8] = 4'h0;
    SS12[6][8] = 4'hC;
    SS12[7][8] = 4'hC;
    SS12[8][8] = 4'hC;
    SS12[9][8] = 4'hC;
    SS12[10][8] = 4'hC;
    SS12[11][8] = 4'hC;
    SS12[12][8] = 4'hC;
    SS12[13][8] = 4'h0;
    SS12[14][8] = 4'hD;
    SS12[15][8] = 4'hD;
    SS12[16][8] = 4'hD;
    SS12[17][8] = 4'h0;
    SS12[18][8] = 4'h0;
    SS12[19][8] = 4'h0;
    SS12[20][8] = 4'h0;
    SS12[21][8] = 4'h0;
    SS12[22][8] = 4'h0;
    SS12[23][8] = 4'h0;
    SS12[24][8] = 4'h0;
    SS12[25][8] = 4'h0;
    SS12[26][8] = 4'h0;
    SS12[27][8] = 4'h0;
    SS12[28][8] = 4'h0;
    SS12[29][8] = 4'h0;
    SS12[30][8] = 4'h0;
    SS12[31][8] = 4'h0;
    SS12[32][8] = 4'h0;
    SS12[33][8] = 4'h0;
    SS12[34][8] = 4'h0;
    SS12[35][8] = 4'h0;
    SS12[36][8] = 4'h0;
    SS12[37][8] = 4'h0;
    SS12[38][8] = 4'h0;
    SS12[39][8] = 4'h0;
    SS12[40][8] = 4'h0;
    SS12[41][8] = 4'h0;
    SS12[42][8] = 4'h0;
    SS12[43][8] = 4'h0;
    SS12[44][8] = 4'h0;
    SS12[45][8] = 4'h0;
    SS12[46][8] = 4'h0;
    SS12[47][8] = 4'h0;
    SS12[0][9] = 4'h0;
    SS12[1][9] = 4'h0;
    SS12[2][9] = 4'h0;
    SS12[3][9] = 4'h0;
    SS12[4][9] = 4'h0;
    SS12[5][9] = 4'hC;
    SS12[6][9] = 4'hC;
    SS12[7][9] = 4'hC;
    SS12[8][9] = 4'hC;
    SS12[9][9] = 4'hC;
    SS12[10][9] = 4'hC;
    SS12[11][9] = 4'hC;
    SS12[12][9] = 4'hC;
    SS12[13][9] = 4'hC;
    SS12[14][9] = 4'hD;
    SS12[15][9] = 4'hD;
    SS12[16][9] = 4'hD;
    SS12[17][9] = 4'hD;
    SS12[18][9] = 4'h0;
    SS12[19][9] = 4'h0;
    SS12[20][9] = 4'h0;
    SS12[21][9] = 4'h0;
    SS12[22][9] = 4'h0;
    SS12[23][9] = 4'h0;
    SS12[24][9] = 4'h0;
    SS12[25][9] = 4'h0;
    SS12[26][9] = 4'h0;
    SS12[27][9] = 4'h0;
    SS12[28][9] = 4'h0;
    SS12[29][9] = 4'h0;
    SS12[30][9] = 4'h0;
    SS12[31][9] = 4'h0;
    SS12[32][9] = 4'h0;
    SS12[33][9] = 4'h0;
    SS12[34][9] = 4'h0;
    SS12[35][9] = 4'h0;
    SS12[36][9] = 4'h0;
    SS12[37][9] = 4'h0;
    SS12[38][9] = 4'h0;
    SS12[39][9] = 4'h0;
    SS12[40][9] = 4'h0;
    SS12[41][9] = 4'h0;
    SS12[42][9] = 4'h0;
    SS12[43][9] = 4'h0;
    SS12[44][9] = 4'h0;
    SS12[45][9] = 4'h0;
    SS12[46][9] = 4'h0;
    SS12[47][9] = 4'h0;
    SS12[0][10] = 4'h0;
    SS12[1][10] = 4'h0;
    SS12[2][10] = 4'h0;
    SS12[3][10] = 4'h0;
    SS12[4][10] = 4'h0;
    SS12[5][10] = 4'h0;
    SS12[6][10] = 4'hC;
    SS12[7][10] = 4'hC;
    SS12[8][10] = 4'hC;
    SS12[9][10] = 4'hC;
    SS12[10][10] = 4'hC;
    SS12[11][10] = 4'hC;
    SS12[12][10] = 4'hC;
    SS12[13][10] = 4'hC;
    SS12[14][10] = 4'hC;
    SS12[15][10] = 4'hD;
    SS12[16][10] = 4'hD;
    SS12[17][10] = 4'hD;
    SS12[18][10] = 4'hD;
    SS12[19][10] = 4'h0;
    SS12[20][10] = 4'h0;
    SS12[21][10] = 4'h0;
    SS12[22][10] = 4'h0;
    SS12[23][10] = 4'h0;
    SS12[24][10] = 4'h0;
    SS12[25][10] = 4'h0;
    SS12[26][10] = 4'h0;
    SS12[27][10] = 4'h0;
    SS12[28][10] = 4'h0;
    SS12[29][10] = 4'h0;
    SS12[30][10] = 4'h0;
    SS12[31][10] = 4'h0;
    SS12[32][10] = 4'h0;
    SS12[33][10] = 4'h0;
    SS12[34][10] = 4'h0;
    SS12[35][10] = 4'h0;
    SS12[36][10] = 4'h0;
    SS12[37][10] = 4'h0;
    SS12[38][10] = 4'h0;
    SS12[39][10] = 4'h0;
    SS12[40][10] = 4'h0;
    SS12[41][10] = 4'h0;
    SS12[42][10] = 4'h0;
    SS12[43][10] = 4'h0;
    SS12[44][10] = 4'h0;
    SS12[45][10] = 4'h0;
    SS12[46][10] = 4'h0;
    SS12[47][10] = 4'h0;
    SS12[0][11] = 4'h0;
    SS12[1][11] = 4'h0;
    SS12[2][11] = 4'h0;
    SS12[3][11] = 4'h0;
    SS12[4][11] = 4'h0;
    SS12[5][11] = 4'h0;
    SS12[6][11] = 4'h0;
    SS12[7][11] = 4'hC;
    SS12[8][11] = 4'hC;
    SS12[9][11] = 4'hC;
    SS12[10][11] = 4'hC;
    SS12[11][11] = 4'hC;
    SS12[12][11] = 4'hC;
    SS12[13][11] = 4'hC;
    SS12[14][11] = 4'hC;
    SS12[15][11] = 4'hC;
    SS12[16][11] = 4'hD;
    SS12[17][11] = 4'hD;
    SS12[18][11] = 4'hD;
    SS12[19][11] = 4'hD;
    SS12[20][11] = 4'h0;
    SS12[21][11] = 4'h0;
    SS12[22][11] = 4'h0;
    SS12[23][11] = 4'h0;
    SS12[24][11] = 4'h0;
    SS12[25][11] = 4'h0;
    SS12[26][11] = 4'h0;
    SS12[27][11] = 4'h0;
    SS12[28][11] = 4'h2;
    SS12[29][11] = 4'h0;
    SS12[30][11] = 4'h0;
    SS12[31][11] = 4'h0;
    SS12[32][11] = 4'h0;
    SS12[33][11] = 4'h0;
    SS12[34][11] = 4'h0;
    SS12[35][11] = 4'h0;
    SS12[36][11] = 4'h2;
    SS12[37][11] = 4'h0;
    SS12[38][11] = 4'h0;
    SS12[39][11] = 4'h0;
    SS12[40][11] = 4'h0;
    SS12[41][11] = 4'h0;
    SS12[42][11] = 4'h0;
    SS12[43][11] = 4'h0;
    SS12[44][11] = 4'h0;
    SS12[45][11] = 4'h0;
    SS12[46][11] = 4'h0;
    SS12[47][11] = 4'h0;
    SS12[0][12] = 4'h0;
    SS12[1][12] = 4'h0;
    SS12[2][12] = 4'h0;
    SS12[3][12] = 4'h0;
    SS12[4][12] = 4'h0;
    SS12[5][12] = 4'h0;
    SS12[6][12] = 4'h0;
    SS12[7][12] = 4'h0;
    SS12[8][12] = 4'hC;
    SS12[9][12] = 4'hC;
    SS12[10][12] = 4'hC;
    SS12[11][12] = 4'hC;
    SS12[12][12] = 4'hC;
    SS12[13][12] = 4'hC;
    SS12[14][12] = 4'hC;
    SS12[15][12] = 4'hC;
    SS12[16][12] = 4'hC;
    SS12[17][12] = 4'hD;
    SS12[18][12] = 4'hD;
    SS12[19][12] = 4'hD;
    SS12[20][12] = 4'hD;
    SS12[21][12] = 4'h0;
    SS12[22][12] = 4'h0;
    SS12[23][12] = 4'h0;
    SS12[24][12] = 4'h0;
    SS12[25][12] = 4'h0;
    SS12[26][12] = 4'h0;
    SS12[27][12] = 4'h3;
    SS12[28][12] = 4'h3;
    SS12[29][12] = 4'h2;
    SS12[30][12] = 4'h0;
    SS12[31][12] = 4'h0;
    SS12[32][12] = 4'h0;
    SS12[33][12] = 4'h0;
    SS12[34][12] = 4'h0;
    SS12[35][12] = 4'h2;
    SS12[36][12] = 4'h3;
    SS12[37][12] = 4'h3;
    SS12[38][12] = 4'h0;
    SS12[39][12] = 4'h0;
    SS12[40][12] = 4'hD;
    SS12[41][12] = 4'hD;
    SS12[42][12] = 4'h0;
    SS12[43][12] = 4'h0;
    SS12[44][12] = 4'hD;
    SS12[45][12] = 4'hD;
    SS12[46][12] = 4'h0;
    SS12[47][12] = 4'h0;
    SS12[0][13] = 4'h0;
    SS12[1][13] = 4'h0;
    SS12[2][13] = 4'h0;
    SS12[3][13] = 4'h0;
    SS12[4][13] = 4'h0;
    SS12[5][13] = 4'h0;
    SS12[6][13] = 4'h0;
    SS12[7][13] = 4'h0;
    SS12[8][13] = 4'h0;
    SS12[9][13] = 4'hC;
    SS12[10][13] = 4'hC;
    SS12[11][13] = 4'hC;
    SS12[12][13] = 4'hC;
    SS12[13][13] = 4'hC;
    SS12[14][13] = 4'hC;
    SS12[15][13] = 4'hC;
    SS12[16][13] = 4'hC;
    SS12[17][13] = 4'hC;
    SS12[18][13] = 4'hD;
    SS12[19][13] = 4'hD;
    SS12[20][13] = 4'hD;
    SS12[21][13] = 4'hD;
    SS12[22][13] = 4'h0;
    SS12[23][13] = 4'h0;
    SS12[24][13] = 4'h0;
    SS12[25][13] = 4'h0;
    SS12[26][13] = 4'h3;
    SS12[27][13] = 4'h3;
    SS12[28][13] = 4'h3;
    SS12[29][13] = 4'h3;
    SS12[30][13] = 4'h0;
    SS12[31][13] = 4'h0;
    SS12[32][13] = 4'h0;
    SS12[33][13] = 4'h0;
    SS12[34][13] = 4'hE;
    SS12[35][13] = 4'h3;
    SS12[36][13] = 4'h3;
    SS12[37][13] = 4'h3;
    SS12[38][13] = 4'h3;
    SS12[39][13] = 4'hD;
    SS12[40][13] = 4'hD;
    SS12[41][13] = 4'hD;
    SS12[42][13] = 4'hD;
    SS12[43][13] = 4'hD;
    SS12[44][13] = 4'hD;
    SS12[45][13] = 4'hD;
    SS12[46][13] = 4'hD;
    SS12[47][13] = 4'h0;
    SS12[0][14] = 4'h0;
    SS12[1][14] = 4'h0;
    SS12[2][14] = 4'h0;
    SS12[3][14] = 4'h0;
    SS12[4][14] = 4'h0;
    SS12[5][14] = 4'h0;
    SS12[6][14] = 4'h0;
    SS12[7][14] = 4'h0;
    SS12[8][14] = 4'hD;
    SS12[9][14] = 4'hD;
    SS12[10][14] = 4'hC;
    SS12[11][14] = 4'hC;
    SS12[12][14] = 4'hC;
    SS12[13][14] = 4'hC;
    SS12[14][14] = 4'hC;
    SS12[15][14] = 4'hC;
    SS12[16][14] = 4'hC;
    SS12[17][14] = 4'hC;
    SS12[18][14] = 4'hC;
    SS12[19][14] = 4'hD;
    SS12[20][14] = 4'hD;
    SS12[21][14] = 4'hC;
    SS12[22][14] = 4'hC;
    SS12[23][14] = 4'h0;
    SS12[24][14] = 4'h0;
    SS12[25][14] = 4'hD;
    SS12[26][14] = 4'hD;
    SS12[27][14] = 4'h3;
    SS12[28][14] = 4'h3;
    SS12[29][14] = 4'hD;
    SS12[30][14] = 4'hD;
    SS12[31][14] = 4'h0;
    SS12[32][14] = 4'h0;
    SS12[33][14] = 4'hE;
    SS12[34][14] = 4'hD;
    SS12[35][14] = 4'hD;
    SS12[36][14] = 4'h3;
    SS12[37][14] = 4'h3;
    SS12[38][14] = 4'hD;
    SS12[39][14] = 4'hD;
    SS12[40][14] = 4'hD;
    SS12[41][14] = 4'hD;
    SS12[42][14] = 4'hD;
    SS12[43][14] = 4'hD;
    SS12[44][14] = 4'hD;
    SS12[45][14] = 4'hD;
    SS12[46][14] = 4'h0;
    SS12[47][14] = 4'h0;
    SS12[0][15] = 4'h0;
    SS12[1][15] = 4'h0;
    SS12[2][15] = 4'h0;
    SS12[3][15] = 4'h0;
    SS12[4][15] = 4'h0;
    SS12[5][15] = 4'h0;
    SS12[6][15] = 4'h0;
    SS12[7][15] = 4'hD;
    SS12[8][15] = 4'hD;
    SS12[9][15] = 4'hD;
    SS12[10][15] = 4'hD;
    SS12[11][15] = 4'hC;
    SS12[12][15] = 4'hC;
    SS12[13][15] = 4'hC;
    SS12[14][15] = 4'hC;
    SS12[15][15] = 4'hC;
    SS12[16][15] = 4'hC;
    SS12[17][15] = 4'hC;
    SS12[18][15] = 4'hC;
    SS12[19][15] = 4'hC;
    SS12[20][15] = 4'hC;
    SS12[21][15] = 4'hC;
    SS12[22][15] = 4'hC;
    SS12[23][15] = 4'hC;
    SS12[24][15] = 4'hD;
    SS12[25][15] = 4'hD;
    SS12[26][15] = 4'hD;
    SS12[27][15] = 4'hD;
    SS12[28][15] = 4'hD;
    SS12[29][15] = 4'hD;
    SS12[30][15] = 4'hD;
    SS12[31][15] = 4'hD;
    SS12[32][15] = 4'hD;
    SS12[33][15] = 4'hD;
    SS12[34][15] = 4'hD;
    SS12[35][15] = 4'hD;
    SS12[36][15] = 4'hD;
    SS12[37][15] = 4'hD;
    SS12[38][15] = 4'hD;
    SS12[39][15] = 4'hD;
    SS12[40][15] = 4'hD;
    SS12[41][15] = 4'hD;
    SS12[42][15] = 4'hD;
    SS12[43][15] = 4'hD;
    SS12[44][15] = 4'hD;
    SS12[45][15] = 4'h0;
    SS12[46][15] = 4'h0;
    SS12[47][15] = 4'h0;
    SS12[0][16] = 4'h0;
    SS12[1][16] = 4'h0;
    SS12[2][16] = 4'h0;
    SS12[3][16] = 4'h0;
    SS12[4][16] = 4'h0;
    SS12[5][16] = 4'h0;
    SS12[6][16] = 4'h0;
    SS12[7][16] = 4'h0;
    SS12[8][16] = 4'hD;
    SS12[9][16] = 4'hD;
    SS12[10][16] = 4'hD;
    SS12[11][16] = 4'hD;
    SS12[12][16] = 4'hC;
    SS12[13][16] = 4'hC;
    SS12[14][16] = 4'hC;
    SS12[15][16] = 4'hC;
    SS12[16][16] = 4'hC;
    SS12[17][16] = 4'hC;
    SS12[18][16] = 4'hC;
    SS12[19][16] = 4'hC;
    SS12[20][16] = 4'hC;
    SS12[21][16] = 4'hC;
    SS12[22][16] = 4'hC;
    SS12[23][16] = 4'hD;
    SS12[24][16] = 4'hD;
    SS12[25][16] = 4'hD;
    SS12[26][16] = 4'hD;
    SS12[27][16] = 4'hD;
    SS12[28][16] = 4'hD;
    SS12[29][16] = 4'hD;
    SS12[30][16] = 4'hD;
    SS12[31][16] = 4'hD;
    SS12[32][16] = 4'hD;
    SS12[33][16] = 4'hD;
    SS12[34][16] = 4'hD;
    SS12[35][16] = 4'hD;
    SS12[36][16] = 4'hE;
    SS12[37][16] = 4'hE;
    SS12[38][16] = 4'hD;
    SS12[39][16] = 4'hD;
    SS12[40][16] = 4'hE;
    SS12[41][16] = 4'hE;
    SS12[42][16] = 4'hD;
    SS12[43][16] = 4'hD;
    SS12[44][16] = 4'h0;
    SS12[45][16] = 4'h0;
    SS12[46][16] = 4'h0;
    SS12[47][16] = 4'h0;
    SS12[0][17] = 4'h0;
    SS12[1][17] = 4'h0;
    SS12[2][17] = 4'h0;
    SS12[3][17] = 4'h0;
    SS12[4][17] = 4'h0;
    SS12[5][17] = 4'h0;
    SS12[6][17] = 4'h0;
    SS12[7][17] = 4'h0;
    SS12[8][17] = 4'h0;
    SS12[9][17] = 4'hD;
    SS12[10][17] = 4'hD;
    SS12[11][17] = 4'hD;
    SS12[12][17] = 4'hD;
    SS12[13][17] = 4'hC;
    SS12[14][17] = 4'hC;
    SS12[15][17] = 4'hC;
    SS12[16][17] = 4'hC;
    SS12[17][17] = 4'hC;
    SS12[18][17] = 4'hC;
    SS12[19][17] = 4'hC;
    SS12[20][17] = 4'hC;
    SS12[21][17] = 4'hC;
    SS12[22][17] = 4'hD;
    SS12[23][17] = 4'hD;
    SS12[24][17] = 4'hD;
    SS12[25][17] = 4'hD;
    SS12[26][17] = 4'hD;
    SS12[27][17] = 4'hD;
    SS12[28][17] = 4'hD;
    SS12[29][17] = 4'hD;
    SS12[30][17] = 4'hD;
    SS12[31][17] = 4'hD;
    SS12[32][17] = 4'hD;
    SS12[33][17] = 4'hD;
    SS12[34][17] = 4'hD;
    SS12[35][17] = 4'hE;
    SS12[36][17] = 4'hE;
    SS12[37][17] = 4'hE;
    SS12[38][17] = 4'hE;
    SS12[39][17] = 4'hE;
    SS12[40][17] = 4'hE;
    SS12[41][17] = 4'hE;
    SS12[42][17] = 4'hE;
    SS12[43][17] = 4'h0;
    SS12[44][17] = 4'h0;
    SS12[45][17] = 4'h0;
    SS12[46][17] = 4'h0;
    SS12[47][17] = 4'h0;
    SS12[0][18] = 4'h0;
    SS12[1][18] = 4'h0;
    SS12[2][18] = 4'h0;
    SS12[3][18] = 4'h0;
    SS12[4][18] = 4'h0;
    SS12[5][18] = 4'h0;
    SS12[6][18] = 4'h0;
    SS12[7][18] = 4'h0;
    SS12[8][18] = 4'h0;
    SS12[9][18] = 4'h0;
    SS12[10][18] = 4'hD;
    SS12[11][18] = 4'hD;
    SS12[12][18] = 4'hD;
    SS12[13][18] = 4'hD;
    SS12[14][18] = 4'hC;
    SS12[15][18] = 4'hC;
    SS12[16][18] = 4'hC;
    SS12[17][18] = 4'hC;
    SS12[18][18] = 4'hC;
    SS12[19][18] = 4'hC;
    SS12[20][18] = 4'hC;
    SS12[21][18] = 4'hA;
    SS12[22][18] = 4'hA;
    SS12[23][18] = 4'hD;
    SS12[24][18] = 4'hD;
    SS12[25][18] = 4'hC;
    SS12[26][18] = 4'hC;
    SS12[27][18] = 4'hD;
    SS12[28][18] = 4'hD;
    SS12[29][18] = 4'hD;
    SS12[30][18] = 4'hE;
    SS12[31][18] = 4'hD;
    SS12[32][18] = 4'hD;
    SS12[33][18] = 4'hD;
    SS12[34][18] = 4'hE;
    SS12[35][18] = 4'hE;
    SS12[36][18] = 4'hE;
    SS12[37][18] = 4'hE;
    SS12[38][18] = 4'hE;
    SS12[39][18] = 4'hE;
    SS12[40][18] = 4'hE;
    SS12[41][18] = 4'hE;
    SS12[42][18] = 4'h0;
    SS12[43][18] = 4'h0;
    SS12[44][18] = 4'h0;
    SS12[45][18] = 4'h0;
    SS12[46][18] = 4'h0;
    SS12[47][18] = 4'h0;
    SS12[0][19] = 4'h0;
    SS12[1][19] = 4'h0;
    SS12[2][19] = 4'h0;
    SS12[3][19] = 4'h0;
    SS12[4][19] = 4'h0;
    SS12[5][19] = 4'h0;
    SS12[6][19] = 4'h0;
    SS12[7][19] = 4'h0;
    SS12[8][19] = 4'h0;
    SS12[9][19] = 4'h0;
    SS12[10][19] = 4'h0;
    SS12[11][19] = 4'hD;
    SS12[12][19] = 4'hD;
    SS12[13][19] = 4'hD;
    SS12[14][19] = 4'hD;
    SS12[15][19] = 4'hC;
    SS12[16][19] = 4'hC;
    SS12[17][19] = 4'hC;
    SS12[18][19] = 4'hC;
    SS12[19][19] = 4'hC;
    SS12[20][19] = 4'hA;
    SS12[21][19] = 4'hA;
    SS12[22][19] = 4'hA;
    SS12[23][19] = 4'hA;
    SS12[24][19] = 4'hC;
    SS12[25][19] = 4'hC;
    SS12[26][19] = 4'hC;
    SS12[27][19] = 4'hC;
    SS12[28][19] = 4'hD;
    SS12[29][19] = 4'hE;
    SS12[30][19] = 4'hE;
    SS12[31][19] = 4'hE;
    SS12[32][19] = 4'hD;
    SS12[33][19] = 4'hE;
    SS12[34][19] = 4'hE;
    SS12[35][19] = 4'hE;
    SS12[36][19] = 4'hE;
    SS12[37][19] = 4'hE;
    SS12[38][19] = 4'hE;
    SS12[39][19] = 4'hE;
    SS12[40][19] = 4'hE;
    SS12[41][19] = 4'h0;
    SS12[42][19] = 4'h0;
    SS12[43][19] = 4'h0;
    SS12[44][19] = 4'h0;
    SS12[45][19] = 4'h0;
    SS12[46][19] = 4'h0;
    SS12[47][19] = 4'h0;
    SS12[0][20] = 4'h0;
    SS12[1][20] = 4'h0;
    SS12[2][20] = 4'h0;
    SS12[3][20] = 4'h0;
    SS12[4][20] = 4'h0;
    SS12[5][20] = 4'h0;
    SS12[6][20] = 4'h0;
    SS12[7][20] = 4'h0;
    SS12[8][20] = 4'h0;
    SS12[9][20] = 4'h0;
    SS12[10][20] = 4'h0;
    SS12[11][20] = 4'h0;
    SS12[12][20] = 4'hD;
    SS12[13][20] = 4'hD;
    SS12[14][20] = 4'hD;
    SS12[15][20] = 4'hC;
    SS12[16][20] = 4'hC;
    SS12[17][20] = 4'hC;
    SS12[18][20] = 4'hC;
    SS12[19][20] = 4'hA;
    SS12[20][20] = 4'hA;
    SS12[21][20] = 4'hA;
    SS12[22][20] = 4'hA;
    SS12[23][20] = 4'hD;
    SS12[24][20] = 4'hD;
    SS12[25][20] = 4'hC;
    SS12[26][20] = 4'hC;
    SS12[27][20] = 4'hC;
    SS12[28][20] = 4'hC;
    SS12[29][20] = 4'hE;
    SS12[30][20] = 4'hE;
    SS12[31][20] = 4'hE;
    SS12[32][20] = 4'hC;
    SS12[33][20] = 4'hE;
    SS12[34][20] = 4'hE;
    SS12[35][20] = 4'hE;
    SS12[36][20] = 4'hC;
    SS12[37][20] = 4'hE;
    SS12[38][20] = 4'hE;
    SS12[39][20] = 4'hE;
    SS12[40][20] = 4'h0;
    SS12[41][20] = 4'h0;
    SS12[42][20] = 4'h0;
    SS12[43][20] = 4'h0;
    SS12[44][20] = 4'h0;
    SS12[45][20] = 4'h0;
    SS12[46][20] = 4'h0;
    SS12[47][20] = 4'h0;
    SS12[0][21] = 4'h0;
    SS12[1][21] = 4'h0;
    SS12[2][21] = 4'h0;
    SS12[3][21] = 4'h0;
    SS12[4][21] = 4'h0;
    SS12[5][21] = 4'h0;
    SS12[6][21] = 4'h0;
    SS12[7][21] = 4'h0;
    SS12[8][21] = 4'h0;
    SS12[9][21] = 4'h0;
    SS12[10][21] = 4'h0;
    SS12[11][21] = 4'h0;
    SS12[12][21] = 4'h0;
    SS12[13][21] = 4'hD;
    SS12[14][21] = 4'hC;
    SS12[15][21] = 4'hC;
    SS12[16][21] = 4'hC;
    SS12[17][21] = 4'hC;
    SS12[18][21] = 4'hA;
    SS12[19][21] = 4'hA;
    SS12[20][21] = 4'hA;
    SS12[21][21] = 4'hA;
    SS12[22][21] = 4'hD;
    SS12[23][21] = 4'hD;
    SS12[24][21] = 4'hD;
    SS12[25][21] = 4'hD;
    SS12[26][21] = 4'hC;
    SS12[27][21] = 4'hC;
    SS12[28][21] = 4'hC;
    SS12[29][21] = 4'hC;
    SS12[30][21] = 4'hE;
    SS12[31][21] = 4'hC;
    SS12[32][21] = 4'hC;
    SS12[33][21] = 4'hC;
    SS12[34][21] = 4'hE;
    SS12[35][21] = 4'hC;
    SS12[36][21] = 4'hC;
    SS12[37][21] = 4'hC;
    SS12[38][21] = 4'hE;
    SS12[39][21] = 4'h0;
    SS12[40][21] = 4'h0;
    SS12[41][21] = 4'h0;
    SS12[42][21] = 4'h0;
    SS12[43][21] = 4'h0;
    SS12[44][21] = 4'h0;
    SS12[45][21] = 4'h0;
    SS12[46][21] = 4'h0;
    SS12[47][21] = 4'h0;
    SS12[0][22] = 4'h0;
    SS12[1][22] = 4'h0;
    SS12[2][22] = 4'h0;
    SS12[3][22] = 4'h0;
    SS12[4][22] = 4'h0;
    SS12[5][22] = 4'h0;
    SS12[6][22] = 4'h0;
    SS12[7][22] = 4'h0;
    SS12[8][22] = 4'h0;
    SS12[9][22] = 4'h0;
    SS12[10][22] = 4'h0;
    SS12[11][22] = 4'h0;
    SS12[12][22] = 4'h0;
    SS12[13][22] = 4'h0;
    SS12[14][22] = 4'hC;
    SS12[15][22] = 4'hC;
    SS12[16][22] = 4'hC;
    SS12[17][22] = 4'hD;
    SS12[18][22] = 4'hA;
    SS12[19][22] = 4'hA;
    SS12[20][22] = 4'hA;
    SS12[21][22] = 4'hD;
    SS12[22][22] = 4'hD;
    SS12[23][22] = 4'hD;
    SS12[24][22] = 4'hD;
    SS12[25][22] = 4'hC;
    SS12[26][22] = 4'hC;
    SS12[27][22] = 4'hC;
    SS12[28][22] = 4'hC;
    SS12[29][22] = 4'hC;
    SS12[30][22] = 4'hC;
    SS12[31][22] = 4'hC;
    SS12[32][22] = 4'hC;
    SS12[33][22] = 4'hC;
    SS12[34][22] = 4'hC;
    SS12[35][22] = 4'hC;
    SS12[36][22] = 4'hC;
    SS12[37][22] = 4'hC;
    SS12[38][22] = 4'hC;
    SS12[39][22] = 4'hD;
    SS12[40][22] = 4'h0;
    SS12[41][22] = 4'h0;
    SS12[42][22] = 4'h0;
    SS12[43][22] = 4'h0;
    SS12[44][22] = 4'h0;
    SS12[45][22] = 4'h0;
    SS12[46][22] = 4'h0;
    SS12[47][22] = 4'h0;
    SS12[0][23] = 4'h0;
    SS12[1][23] = 4'h0;
    SS12[2][23] = 4'h0;
    SS12[3][23] = 4'h0;
    SS12[4][23] = 4'h0;
    SS12[5][23] = 4'h0;
    SS12[6][23] = 4'h0;
    SS12[7][23] = 4'h0;
    SS12[8][23] = 4'h0;
    SS12[9][23] = 4'h0;
    SS12[10][23] = 4'h0;
    SS12[11][23] = 4'h0;
    SS12[12][23] = 4'h0;
    SS12[13][23] = 4'h0;
    SS12[14][23] = 4'h0;
    SS12[15][23] = 4'hC;
    SS12[16][23] = 4'hD;
    SS12[17][23] = 4'hD;
    SS12[18][23] = 4'hD;
    SS12[19][23] = 4'hA;
    SS12[20][23] = 4'hD;
    SS12[21][23] = 4'hD;
    SS12[22][23] = 4'hD;
    SS12[23][23] = 4'hD;
    SS12[24][23] = 4'hC;
    SS12[25][23] = 4'hC;
    SS12[26][23] = 4'hC;
    SS12[27][23] = 4'hC;
    SS12[28][23] = 4'hC;
    SS12[29][23] = 4'hC;
    SS12[30][23] = 4'hC;
    SS12[31][23] = 4'hC;
    SS12[32][23] = 4'hC;
    SS12[33][23] = 4'hC;
    SS12[34][23] = 4'hC;
    SS12[35][23] = 4'hC;
    SS12[36][23] = 4'hC;
    SS12[37][23] = 4'hC;
    SS12[38][23] = 4'hC;
    SS12[39][23] = 4'hC;
    SS12[40][23] = 4'hD;
    SS12[41][23] = 4'h0;
    SS12[42][23] = 4'h0;
    SS12[43][23] = 4'h0;
    SS12[44][23] = 4'h0;
    SS12[45][23] = 4'h0;
    SS12[46][23] = 4'h0;
    SS12[47][23] = 4'h0;
    SS12[0][24] = 4'h0;
    SS12[1][24] = 4'h0;
    SS12[2][24] = 4'h0;
    SS12[3][24] = 4'h0;
    SS12[4][24] = 4'h0;
    SS12[5][24] = 4'h0;
    SS12[6][24] = 4'h0;
    SS12[7][24] = 4'h0;
    SS12[8][24] = 4'h0;
    SS12[9][24] = 4'h0;
    SS12[10][24] = 4'h0;
    SS12[11][24] = 4'h0;
    SS12[12][24] = 4'h0;
    SS12[13][24] = 4'h0;
    SS12[14][24] = 4'h0;
    SS12[15][24] = 4'hD;
    SS12[16][24] = 4'hD;
    SS12[17][24] = 4'hD;
    SS12[18][24] = 4'hD;
    SS12[19][24] = 4'hC;
    SS12[20][24] = 4'hD;
    SS12[21][24] = 4'hD;
    SS12[22][24] = 4'hD;
    SS12[23][24] = 4'hC;
    SS12[24][24] = 4'hC;
    SS12[25][24] = 4'hC;
    SS12[26][24] = 4'hC;
    SS12[27][24] = 4'hC;
    SS12[28][24] = 4'hD;
    SS12[29][24] = 4'hC;
    SS12[30][24] = 4'hC;
    SS12[31][24] = 4'hC;
    SS12[32][24] = 4'hC;
    SS12[33][24] = 4'hC;
    SS12[34][24] = 4'hC;
    SS12[35][24] = 4'hC;
    SS12[36][24] = 4'hC;
    SS12[37][24] = 4'hC;
    SS12[38][24] = 4'hC;
    SS12[39][24] = 4'hC;
    SS12[40][24] = 4'hC;
    SS12[41][24] = 4'h0;
    SS12[42][24] = 4'h0;
    SS12[43][24] = 4'h0;
    SS12[44][24] = 4'h0;
    SS12[45][24] = 4'hC;
    SS12[46][24] = 4'h0;
    SS12[47][24] = 4'h0;
    SS12[0][25] = 4'h0;
    SS12[1][25] = 4'h0;
    SS12[2][25] = 4'h0;
    SS12[3][25] = 4'h0;
    SS12[4][25] = 4'h0;
    SS12[5][25] = 4'h0;
    SS12[6][25] = 4'h0;
    SS12[7][25] = 4'h0;
    SS12[8][25] = 4'h0;
    SS12[9][25] = 4'h0;
    SS12[10][25] = 4'h0;
    SS12[11][25] = 4'h0;
    SS12[12][25] = 4'h0;
    SS12[13][25] = 4'h0;
    SS12[14][25] = 4'hD;
    SS12[15][25] = 4'hD;
    SS12[16][25] = 4'hD;
    SS12[17][25] = 4'hD;
    SS12[18][25] = 4'hC;
    SS12[19][25] = 4'hC;
    SS12[20][25] = 4'hC;
    SS12[21][25] = 4'hD;
    SS12[22][25] = 4'hC;
    SS12[23][25] = 4'hC;
    SS12[24][25] = 4'hC;
    SS12[25][25] = 4'hC;
    SS12[26][25] = 4'hC;
    SS12[27][25] = 4'hD;
    SS12[28][25] = 4'hD;
    SS12[29][25] = 4'hD;
    SS12[30][25] = 4'hC;
    SS12[31][25] = 4'hC;
    SS12[32][25] = 4'hC;
    SS12[33][25] = 4'hC;
    SS12[34][25] = 4'hC;
    SS12[35][25] = 4'hC;
    SS12[36][25] = 4'hC;
    SS12[37][25] = 4'hC;
    SS12[38][25] = 4'hC;
    SS12[39][25] = 4'hC;
    SS12[40][25] = 4'hC;
    SS12[41][25] = 4'hC;
    SS12[42][25] = 4'h0;
    SS12[43][25] = 4'h0;
    SS12[44][25] = 4'hC;
    SS12[45][25] = 4'hC;
    SS12[46][25] = 4'hC;
    SS12[47][25] = 4'h0;
    SS12[0][26] = 4'h0;
    SS12[1][26] = 4'h0;
    SS12[2][26] = 4'h0;
    SS12[3][26] = 4'h0;
    SS12[4][26] = 4'h0;
    SS12[5][26] = 4'h0;
    SS12[6][26] = 4'h0;
    SS12[7][26] = 4'h0;
    SS12[8][26] = 4'h0;
    SS12[9][26] = 4'h0;
    SS12[10][26] = 4'h0;
    SS12[11][26] = 4'h0;
    SS12[12][26] = 4'h0;
    SS12[13][26] = 4'h3;
    SS12[14][26] = 4'hD;
    SS12[15][26] = 4'hD;
    SS12[16][26] = 4'hD;
    SS12[17][26] = 4'hD;
    SS12[18][26] = 4'hC;
    SS12[19][26] = 4'hC;
    SS12[20][26] = 4'hC;
    SS12[21][26] = 4'hC;
    SS12[22][26] = 4'hC;
    SS12[23][26] = 4'hC;
    SS12[24][26] = 4'hC;
    SS12[25][26] = 4'hC;
    SS12[26][26] = 4'hD;
    SS12[27][26] = 4'hD;
    SS12[28][26] = 4'hD;
    SS12[29][26] = 4'hD;
    SS12[30][26] = 4'hE;
    SS12[31][26] = 4'hC;
    SS12[32][26] = 4'hC;
    SS12[33][26] = 4'hC;
    SS12[34][26] = 4'hD;
    SS12[35][26] = 4'hC;
    SS12[36][26] = 4'hC;
    SS12[37][26] = 4'hC;
    SS12[38][26] = 4'hD;
    SS12[39][26] = 4'hC;
    SS12[40][26] = 4'hC;
    SS12[41][26] = 4'hC;
    SS12[42][26] = 4'hC;
    SS12[43][26] = 4'hC;
    SS12[44][26] = 4'hC;
    SS12[45][26] = 4'hC;
    SS12[46][26] = 4'hC;
    SS12[47][26] = 4'hC;
    SS12[0][27] = 4'h0;
    SS12[1][27] = 4'h0;
    SS12[2][27] = 4'h0;
    SS12[3][27] = 4'h0;
    SS12[4][27] = 4'h0;
    SS12[5][27] = 4'h0;
    SS12[6][27] = 4'h0;
    SS12[7][27] = 4'h0;
    SS12[8][27] = 4'h0;
    SS12[9][27] = 4'h0;
    SS12[10][27] = 4'h0;
    SS12[11][27] = 4'h0;
    SS12[12][27] = 4'h3;
    SS12[13][27] = 4'h3;
    SS12[14][27] = 4'h3;
    SS12[15][27] = 4'hD;
    SS12[16][27] = 4'hD;
    SS12[17][27] = 4'hD;
    SS12[18][27] = 4'hD;
    SS12[19][27] = 4'hC;
    SS12[20][27] = 4'hC;
    SS12[21][27] = 4'hC;
    SS12[22][27] = 4'hC;
    SS12[23][27] = 4'hC;
    SS12[24][27] = 4'hC;
    SS12[25][27] = 4'hD;
    SS12[26][27] = 4'hD;
    SS12[27][27] = 4'hD;
    SS12[28][27] = 4'hD;
    SS12[29][27] = 4'hE;
    SS12[30][27] = 4'hE;
    SS12[31][27] = 4'hE;
    SS12[32][27] = 4'hC;
    SS12[33][27] = 4'hD;
    SS12[34][27] = 4'hD;
    SS12[35][27] = 4'hD;
    SS12[36][27] = 4'hC;
    SS12[37][27] = 4'hD;
    SS12[38][27] = 4'hD;
    SS12[39][27] = 4'hD;
    SS12[40][27] = 4'hC;
    SS12[41][27] = 4'hC;
    SS12[42][27] = 4'hC;
    SS12[43][27] = 4'hC;
    SS12[44][27] = 4'hC;
    SS12[45][27] = 4'hC;
    SS12[46][27] = 4'hC;
    SS12[47][27] = 4'hC;
    SS12[0][28] = 4'h0;
    SS12[1][28] = 4'h0;
    SS12[2][28] = 4'h0;
    SS12[3][28] = 4'h0;
    SS12[4][28] = 4'h0;
    SS12[5][28] = 4'h0;
    SS12[6][28] = 4'h0;
    SS12[7][28] = 4'h0;
    SS12[8][28] = 4'h0;
    SS12[9][28] = 4'h0;
    SS12[10][28] = 4'h0;
    SS12[11][28] = 4'h2;
    SS12[12][28] = 4'h3;
    SS12[13][28] = 4'h3;
    SS12[14][28] = 4'h3;
    SS12[15][28] = 4'hD;
    SS12[16][28] = 4'hD;
    SS12[17][28] = 4'hD;
    SS12[18][28] = 4'hD;
    SS12[19][28] = 4'hD;
    SS12[20][28] = 4'hC;
    SS12[21][28] = 4'hC;
    SS12[22][28] = 4'hC;
    SS12[23][28] = 4'hC;
    SS12[24][28] = 4'hD;
    SS12[25][28] = 4'hD;
    SS12[26][28] = 4'hD;
    SS12[27][28] = 4'hD;
    SS12[28][28] = 4'hE;
    SS12[29][28] = 4'hE;
    SS12[30][28] = 4'hE;
    SS12[31][28] = 4'hE;
    SS12[32][28] = 4'hE;
    SS12[33][28] = 4'hD;
    SS12[34][28] = 4'hD;
    SS12[35][28] = 4'hD;
    SS12[36][28] = 4'hD;
    SS12[37][28] = 4'hD;
    SS12[38][28] = 4'hD;
    SS12[39][28] = 4'hD;
    SS12[40][28] = 4'hD;
    SS12[41][28] = 4'hC;
    SS12[42][28] = 4'hC;
    SS12[43][28] = 4'hC;
    SS12[44][28] = 4'hC;
    SS12[45][28] = 4'hC;
    SS12[46][28] = 4'hC;
    SS12[47][28] = 4'hC;
    SS12[0][29] = 4'h0;
    SS12[1][29] = 4'h0;
    SS12[2][29] = 4'h0;
    SS12[3][29] = 4'h0;
    SS12[4][29] = 4'h0;
    SS12[5][29] = 4'h0;
    SS12[6][29] = 4'h0;
    SS12[7][29] = 4'h0;
    SS12[8][29] = 4'h0;
    SS12[9][29] = 4'h0;
    SS12[10][29] = 4'h0;
    SS12[11][29] = 4'h0;
    SS12[12][29] = 4'h2;
    SS12[13][29] = 4'h3;
    SS12[14][29] = 4'hD;
    SS12[15][29] = 4'hD;
    SS12[16][29] = 4'hD;
    SS12[17][29] = 4'hD;
    SS12[18][29] = 4'hD;
    SS12[19][29] = 4'hE;
    SS12[20][29] = 4'hE;
    SS12[21][29] = 4'hC;
    SS12[22][29] = 4'hC;
    SS12[23][29] = 4'hC;
    SS12[24][29] = 4'hC;
    SS12[25][29] = 4'hD;
    SS12[26][29] = 4'hD;
    SS12[27][29] = 4'hE;
    SS12[28][29] = 4'hE;
    SS12[29][29] = 4'hE;
    SS12[30][29] = 4'hE;
    SS12[31][29] = 4'hE;
    SS12[32][29] = 4'hE;
    SS12[33][29] = 4'hE;
    SS12[34][29] = 4'hD;
    SS12[35][29] = 4'hD;
    SS12[36][29] = 4'hE;
    SS12[37][29] = 4'hE;
    SS12[38][29] = 4'hD;
    SS12[39][29] = 4'hD;
    SS12[40][29] = 4'hE;
    SS12[41][29] = 4'hE;
    SS12[42][29] = 4'hC;
    SS12[43][29] = 4'hC;
    SS12[44][29] = 4'hD;
    SS12[45][29] = 4'hD;
    SS12[46][29] = 4'hC;
    SS12[47][29] = 4'hC;
    SS12[0][30] = 4'h0;
    SS12[1][30] = 4'h0;
    SS12[2][30] = 4'h0;
    SS12[3][30] = 4'h0;
    SS12[4][30] = 4'h0;
    SS12[5][30] = 4'h0;
    SS12[6][30] = 4'h0;
    SS12[7][30] = 4'h0;
    SS12[8][30] = 4'h0;
    SS12[9][30] = 4'h0;
    SS12[10][30] = 4'h0;
    SS12[11][30] = 4'h0;
    SS12[12][30] = 4'h0;
    SS12[13][30] = 4'h0;
    SS12[14][30] = 4'hD;
    SS12[15][30] = 4'hD;
    SS12[16][30] = 4'hD;
    SS12[17][30] = 4'hD;
    SS12[18][30] = 4'hE;
    SS12[19][30] = 4'hE;
    SS12[20][30] = 4'hE;
    SS12[21][30] = 4'hE;
    SS12[22][30] = 4'hC;
    SS12[23][30] = 4'hC;
    SS12[24][30] = 4'hC;
    SS12[25][30] = 4'hC;
    SS12[26][30] = 4'hE;
    SS12[27][30] = 4'hE;
    SS12[28][30] = 4'hE;
    SS12[29][30] = 4'hE;
    SS12[30][30] = 4'hE;
    SS12[31][30] = 4'hE;
    SS12[32][30] = 4'hE;
    SS12[33][30] = 4'hE;
    SS12[34][30] = 4'h0;
    SS12[35][30] = 4'hE;
    SS12[36][30] = 4'hE;
    SS12[37][30] = 4'hE;
    SS12[38][30] = 4'hE;
    SS12[39][30] = 4'hE;
    SS12[40][30] = 4'hE;
    SS12[41][30] = 4'hE;
    SS12[42][30] = 4'hE;
    SS12[43][30] = 4'hD;
    SS12[44][30] = 4'hD;
    SS12[45][30] = 4'hD;
    SS12[46][30] = 4'hD;
    SS12[47][30] = 4'hE;
    SS12[0][31] = 4'h0;
    SS12[1][31] = 4'h0;
    SS12[2][31] = 4'h0;
    SS12[3][31] = 4'h0;
    SS12[4][31] = 4'h0;
    SS12[5][31] = 4'h0;
    SS12[6][31] = 4'h0;
    SS12[7][31] = 4'h0;
    SS12[8][31] = 4'h0;
    SS12[9][31] = 4'h0;
    SS12[10][31] = 4'h0;
    SS12[11][31] = 4'h0;
    SS12[12][31] = 4'h0;
    SS12[13][31] = 4'h0;
    SS12[14][31] = 4'h0;
    SS12[15][31] = 4'hD;
    SS12[16][31] = 4'hD;
    SS12[17][31] = 4'hD;
    SS12[18][31] = 4'hD;
    SS12[19][31] = 4'hE;
    SS12[20][31] = 4'hE;
    SS12[21][31] = 4'hC;
    SS12[22][31] = 4'hC;
    SS12[23][31] = 4'hC;
    SS12[24][31] = 4'hC;
    SS12[25][31] = 4'hC;
    SS12[26][31] = 4'hC;
    SS12[27][31] = 4'hE;
    SS12[28][31] = 4'hE;
    SS12[29][31] = 4'hE;
    SS12[30][31] = 4'hE;
    SS12[31][31] = 4'hE;
    SS12[32][31] = 4'hE;
    SS12[33][31] = 4'h0;
    SS12[34][31] = 4'h0;
    SS12[35][31] = 4'h0;
    SS12[36][31] = 4'hE;
    SS12[37][31] = 4'hE;
    SS12[38][31] = 4'h0;
    SS12[39][31] = 4'h0;
    SS12[40][31] = 4'hE;
    SS12[41][31] = 4'hE;
    SS12[42][31] = 4'h0;
    SS12[43][31] = 4'h0;
    SS12[44][31] = 4'hD;
    SS12[45][31] = 4'hD;
    SS12[46][31] = 4'h0;
    SS12[47][31] = 4'h0;
    SS12[0][32] = 4'h0;
    SS12[1][32] = 4'h0;
    SS12[2][32] = 4'h0;
    SS12[3][32] = 4'h0;
    SS12[4][32] = 4'h0;
    SS12[5][32] = 4'h0;
    SS12[6][32] = 4'h0;
    SS12[7][32] = 4'h0;
    SS12[8][32] = 4'h0;
    SS12[9][32] = 4'h0;
    SS12[10][32] = 4'h0;
    SS12[11][32] = 4'h0;
    SS12[12][32] = 4'h0;
    SS12[13][32] = 4'h0;
    SS12[14][32] = 4'h0;
    SS12[15][32] = 4'hD;
    SS12[16][32] = 4'hD;
    SS12[17][32] = 4'hD;
    SS12[18][32] = 4'hD;
    SS12[19][32] = 4'hD;
    SS12[20][32] = 4'hC;
    SS12[21][32] = 4'hC;
    SS12[22][32] = 4'hC;
    SS12[23][32] = 4'hC;
    SS12[24][32] = 4'hC;
    SS12[25][32] = 4'hC;
    SS12[26][32] = 4'hC;
    SS12[27][32] = 4'hC;
    SS12[28][32] = 4'hE;
    SS12[29][32] = 4'hE;
    SS12[30][32] = 4'hE;
    SS12[31][32] = 4'hE;
    SS12[32][32] = 4'hF;
    SS12[33][32] = 4'h0;
    SS12[34][32] = 4'h0;
    SS12[35][32] = 4'h0;
    SS12[36][32] = 4'h0;
    SS12[37][32] = 4'h0;
    SS12[38][32] = 4'h0;
    SS12[39][32] = 4'h0;
    SS12[40][32] = 4'h0;
    SS12[41][32] = 4'h0;
    SS12[42][32] = 4'h0;
    SS12[43][32] = 4'h0;
    SS12[44][32] = 4'h0;
    SS12[45][32] = 4'h0;
    SS12[46][32] = 4'h0;
    SS12[47][32] = 4'h0;
    SS12[0][33] = 4'h0;
    SS12[1][33] = 4'h0;
    SS12[2][33] = 4'h0;
    SS12[3][33] = 4'h0;
    SS12[4][33] = 4'h0;
    SS12[5][33] = 4'h0;
    SS12[6][33] = 4'h0;
    SS12[7][33] = 4'h0;
    SS12[8][33] = 4'h0;
    SS12[9][33] = 4'h0;
    SS12[10][33] = 4'h0;
    SS12[11][33] = 4'h0;
    SS12[12][33] = 4'h0;
    SS12[13][33] = 4'h0;
    SS12[14][33] = 4'hE;
    SS12[15][33] = 4'hD;
    SS12[16][33] = 4'hD;
    SS12[17][33] = 4'hD;
    SS12[18][33] = 4'hD;
    SS12[19][33] = 4'hE;
    SS12[20][33] = 4'hE;
    SS12[21][33] = 4'hC;
    SS12[22][33] = 4'hC;
    SS12[23][33] = 4'hC;
    SS12[24][33] = 4'hC;
    SS12[25][33] = 4'hC;
    SS12[26][33] = 4'hC;
    SS12[27][33] = 4'hD;
    SS12[28][33] = 4'hD;
    SS12[29][33] = 4'hE;
    SS12[30][33] = 4'hE;
    SS12[31][33] = 4'h0;
    SS12[32][33] = 4'h0;
    SS12[33][33] = 4'h0;
    SS12[34][33] = 4'h0;
    SS12[35][33] = 4'h0;
    SS12[36][33] = 4'h0;
    SS12[37][33] = 4'h0;
    SS12[38][33] = 4'h0;
    SS12[39][33] = 4'h0;
    SS12[40][33] = 4'h0;
    SS12[41][33] = 4'h0;
    SS12[42][33] = 4'h0;
    SS12[43][33] = 4'h0;
    SS12[44][33] = 4'h0;
    SS12[45][33] = 4'h0;
    SS12[46][33] = 4'h0;
    SS12[47][33] = 4'h0;
    SS12[0][34] = 4'h0;
    SS12[1][34] = 4'h0;
    SS12[2][34] = 4'h0;
    SS12[3][34] = 4'h0;
    SS12[4][34] = 4'h0;
    SS12[5][34] = 4'h0;
    SS12[6][34] = 4'h0;
    SS12[7][34] = 4'h0;
    SS12[8][34] = 4'h0;
    SS12[9][34] = 4'h0;
    SS12[10][34] = 4'h0;
    SS12[11][34] = 4'h0;
    SS12[12][34] = 4'h0;
    SS12[13][34] = 4'hE;
    SS12[14][34] = 4'hD;
    SS12[15][34] = 4'hD;
    SS12[16][34] = 4'hD;
    SS12[17][34] = 4'hD;
    SS12[18][34] = 4'hE;
    SS12[19][34] = 4'hE;
    SS12[20][34] = 4'hE;
    SS12[21][34] = 4'hE;
    SS12[22][34] = 4'hC;
    SS12[23][34] = 4'hC;
    SS12[24][34] = 4'hC;
    SS12[25][34] = 4'hC;
    SS12[26][34] = 4'hD;
    SS12[27][34] = 4'hD;
    SS12[28][34] = 4'hD;
    SS12[29][34] = 4'hD;
    SS12[30][34] = 4'h0;
    SS12[31][34] = 4'h0;
    SS12[32][34] = 4'h0;
    SS12[33][34] = 4'h0;
    SS12[34][34] = 4'h0;
    SS12[35][34] = 4'h0;
    SS12[36][34] = 4'h0;
    SS12[37][34] = 4'h0;
    SS12[38][34] = 4'h0;
    SS12[39][34] = 4'h0;
    SS12[40][34] = 4'h0;
    SS12[41][34] = 4'h0;
    SS12[42][34] = 4'h0;
    SS12[43][34] = 4'h0;
    SS12[44][34] = 4'h0;
    SS12[45][34] = 4'h0;
    SS12[46][34] = 4'h0;
    SS12[47][34] = 4'h0;
    SS12[0][35] = 4'h0;
    SS12[1][35] = 4'h0;
    SS12[2][35] = 4'h0;
    SS12[3][35] = 4'h0;
    SS12[4][35] = 4'h0;
    SS12[5][35] = 4'h0;
    SS12[6][35] = 4'h0;
    SS12[7][35] = 4'h0;
    SS12[8][35] = 4'h0;
    SS12[9][35] = 4'h0;
    SS12[10][35] = 4'h0;
    SS12[11][35] = 4'h0;
    SS12[12][35] = 4'h2;
    SS12[13][35] = 4'h3;
    SS12[14][35] = 4'hD;
    SS12[15][35] = 4'hD;
    SS12[16][35] = 4'hD;
    SS12[17][35] = 4'hE;
    SS12[18][35] = 4'hE;
    SS12[19][35] = 4'hE;
    SS12[20][35] = 4'hE;
    SS12[21][35] = 4'hC;
    SS12[22][35] = 4'hC;
    SS12[23][35] = 4'hC;
    SS12[24][35] = 4'hC;
    SS12[25][35] = 4'hC;
    SS12[26][35] = 4'hC;
    SS12[27][35] = 4'hD;
    SS12[28][35] = 4'hD;
    SS12[29][35] = 4'hD;
    SS12[30][35] = 4'hE;
    SS12[31][35] = 4'h0;
    SS12[32][35] = 4'h0;
    SS12[33][35] = 4'h0;
    SS12[34][35] = 4'h0;
    SS12[35][35] = 4'h0;
    SS12[36][35] = 4'h0;
    SS12[37][35] = 4'h0;
    SS12[38][35] = 4'h0;
    SS12[39][35] = 4'h0;
    SS12[40][35] = 4'h0;
    SS12[41][35] = 4'h0;
    SS12[42][35] = 4'h0;
    SS12[43][35] = 4'h0;
    SS12[44][35] = 4'h0;
    SS12[45][35] = 4'h0;
    SS12[46][35] = 4'h0;
    SS12[47][35] = 4'h0;
    SS12[0][36] = 4'h0;
    SS12[1][36] = 4'h0;
    SS12[2][36] = 4'h0;
    SS12[3][36] = 4'h0;
    SS12[4][36] = 4'h0;
    SS12[5][36] = 4'h0;
    SS12[6][36] = 4'h0;
    SS12[7][36] = 4'h0;
    SS12[8][36] = 4'h0;
    SS12[9][36] = 4'h0;
    SS12[10][36] = 4'h0;
    SS12[11][36] = 4'h2;
    SS12[12][36] = 4'h3;
    SS12[13][36] = 4'h3;
    SS12[14][36] = 4'h3;
    SS12[15][36] = 4'hD;
    SS12[16][36] = 4'hE;
    SS12[17][36] = 4'hE;
    SS12[18][36] = 4'hE;
    SS12[19][36] = 4'hE;
    SS12[20][36] = 4'hC;
    SS12[21][36] = 4'hC;
    SS12[22][36] = 4'hC;
    SS12[23][36] = 4'hC;
    SS12[24][36] = 4'hC;
    SS12[25][36] = 4'hC;
    SS12[26][36] = 4'hC;
    SS12[27][36] = 4'hC;
    SS12[28][36] = 4'hD;
    SS12[29][36] = 4'hE;
    SS12[30][36] = 4'hE;
    SS12[31][36] = 4'hE;
    SS12[32][36] = 4'h0;
    SS12[33][36] = 4'h0;
    SS12[34][36] = 4'h0;
    SS12[35][36] = 4'h0;
    SS12[36][36] = 4'h0;
    SS12[37][36] = 4'h0;
    SS12[38][36] = 4'h0;
    SS12[39][36] = 4'h0;
    SS12[40][36] = 4'h0;
    SS12[41][36] = 4'h0;
    SS12[42][36] = 4'h0;
    SS12[43][36] = 4'h0;
    SS12[44][36] = 4'h0;
    SS12[45][36] = 4'h0;
    SS12[46][36] = 4'h0;
    SS12[47][36] = 4'h0;
    SS12[0][37] = 4'h0;
    SS12[1][37] = 4'h0;
    SS12[2][37] = 4'h0;
    SS12[3][37] = 4'h0;
    SS12[4][37] = 4'h0;
    SS12[5][37] = 4'h0;
    SS12[6][37] = 4'h0;
    SS12[7][37] = 4'h0;
    SS12[8][37] = 4'h0;
    SS12[9][37] = 4'h0;
    SS12[10][37] = 4'h0;
    SS12[11][37] = 4'h0;
    SS12[12][37] = 4'h3;
    SS12[13][37] = 4'h3;
    SS12[14][37] = 4'h3;
    SS12[15][37] = 4'hD;
    SS12[16][37] = 4'hE;
    SS12[17][37] = 4'hE;
    SS12[18][37] = 4'hE;
    SS12[19][37] = 4'hE;
    SS12[20][37] = 4'hE;
    SS12[21][37] = 4'hC;
    SS12[22][37] = 4'hC;
    SS12[23][37] = 4'hC;
    SS12[24][37] = 4'hC;
    SS12[25][37] = 4'hC;
    SS12[26][37] = 4'hC;
    SS12[27][37] = 4'hD;
    SS12[28][37] = 4'hD;
    SS12[29][37] = 4'hE;
    SS12[30][37] = 4'hE;
    SS12[31][37] = 4'hE;
    SS12[32][37] = 4'h0;
    SS12[33][37] = 4'h0;
    SS12[34][37] = 4'h0;
    SS12[35][37] = 4'h0;
    SS12[36][37] = 4'h0;
    SS12[37][37] = 4'h0;
    SS12[38][37] = 4'h0;
    SS12[39][37] = 4'h0;
    SS12[40][37] = 4'h0;
    SS12[41][37] = 4'h0;
    SS12[42][37] = 4'h0;
    SS12[43][37] = 4'h0;
    SS12[44][37] = 4'h0;
    SS12[45][37] = 4'h0;
    SS12[46][37] = 4'h0;
    SS12[47][37] = 4'h0;
    SS12[0][38] = 4'h0;
    SS12[1][38] = 4'h0;
    SS12[2][38] = 4'h0;
    SS12[3][38] = 4'h0;
    SS12[4][38] = 4'h0;
    SS12[5][38] = 4'h0;
    SS12[6][38] = 4'h0;
    SS12[7][38] = 4'h0;
    SS12[8][38] = 4'h0;
    SS12[9][38] = 4'h0;
    SS12[10][38] = 4'h0;
    SS12[11][38] = 4'h0;
    SS12[12][38] = 4'h0;
    SS12[13][38] = 4'h3;
    SS12[14][38] = 4'hD;
    SS12[15][38] = 4'hD;
    SS12[16][38] = 4'hD;
    SS12[17][38] = 4'hE;
    SS12[18][38] = 4'hE;
    SS12[19][38] = 4'hE;
    SS12[20][38] = 4'hE;
    SS12[21][38] = 4'hE;
    SS12[22][38] = 4'hC;
    SS12[23][38] = 4'hC;
    SS12[24][38] = 4'hC;
    SS12[25][38] = 4'hC;
    SS12[26][38] = 4'hD;
    SS12[27][38] = 4'hD;
    SS12[28][38] = 4'hD;
    SS12[29][38] = 4'hD;
    SS12[30][38] = 4'hE;
    SS12[31][38] = 4'h0;
    SS12[32][38] = 4'h0;
    SS12[33][38] = 4'h0;
    SS12[34][38] = 4'h0;
    SS12[35][38] = 4'h0;
    SS12[36][38] = 4'h0;
    SS12[37][38] = 4'h0;
    SS12[38][38] = 4'h0;
    SS12[39][38] = 4'h0;
    SS12[40][38] = 4'h0;
    SS12[41][38] = 4'h0;
    SS12[42][38] = 4'h0;
    SS12[43][38] = 4'h0;
    SS12[44][38] = 4'h0;
    SS12[45][38] = 4'h0;
    SS12[46][38] = 4'h0;
    SS12[47][38] = 4'h0;
    SS12[0][39] = 4'h0;
    SS12[1][39] = 4'h0;
    SS12[2][39] = 4'h0;
    SS12[3][39] = 4'h0;
    SS12[4][39] = 4'h0;
    SS12[5][39] = 4'h0;
    SS12[6][39] = 4'h0;
    SS12[7][39] = 4'h0;
    SS12[8][39] = 4'h0;
    SS12[9][39] = 4'h0;
    SS12[10][39] = 4'h0;
    SS12[11][39] = 4'h0;
    SS12[12][39] = 4'h0;
    SS12[13][39] = 4'hD;
    SS12[14][39] = 4'hD;
    SS12[15][39] = 4'hD;
    SS12[16][39] = 4'hD;
    SS12[17][39] = 4'hE;
    SS12[18][39] = 4'hE;
    SS12[19][39] = 4'hE;
    SS12[20][39] = 4'hE;
    SS12[21][39] = 4'h0;
    SS12[22][39] = 4'hD;
    SS12[23][39] = 4'hC;
    SS12[24][39] = 4'hC;
    SS12[25][39] = 4'hC;
    SS12[26][39] = 4'hC;
    SS12[27][39] = 4'hD;
    SS12[28][39] = 4'hD;
    SS12[29][39] = 4'hD;
    SS12[30][39] = 4'hE;
    SS12[31][39] = 4'h0;
    SS12[32][39] = 4'h0;
    SS12[33][39] = 4'h0;
    SS12[34][39] = 4'h0;
    SS12[35][39] = 4'h0;
    SS12[36][39] = 4'h0;
    SS12[37][39] = 4'h0;
    SS12[38][39] = 4'h0;
    SS12[39][39] = 4'h0;
    SS12[40][39] = 4'h0;
    SS12[41][39] = 4'h0;
    SS12[42][39] = 4'h0;
    SS12[43][39] = 4'h0;
    SS12[44][39] = 4'h0;
    SS12[45][39] = 4'h0;
    SS12[46][39] = 4'h0;
    SS12[47][39] = 4'h0;
    SS12[0][40] = 4'h0;
    SS12[1][40] = 4'h0;
    SS12[2][40] = 4'h0;
    SS12[3][40] = 4'h0;
    SS12[4][40] = 4'h0;
    SS12[5][40] = 4'h0;
    SS12[6][40] = 4'h0;
    SS12[7][40] = 4'h0;
    SS12[8][40] = 4'h0;
    SS12[9][40] = 4'h0;
    SS12[10][40] = 4'h0;
    SS12[11][40] = 4'h0;
    SS12[12][40] = 4'hD;
    SS12[13][40] = 4'hD;
    SS12[14][40] = 4'hD;
    SS12[15][40] = 4'hD;
    SS12[16][40] = 4'hE;
    SS12[17][40] = 4'hE;
    SS12[18][40] = 4'hE;
    SS12[19][40] = 4'hE;
    SS12[20][40] = 4'h0;
    SS12[21][40] = 4'h0;
    SS12[22][40] = 4'h0;
    SS12[23][40] = 4'hD;
    SS12[24][40] = 4'hC;
    SS12[25][40] = 4'hC;
    SS12[26][40] = 4'hC;
    SS12[27][40] = 4'hC;
    SS12[28][40] = 4'hD;
    SS12[29][40] = 4'hE;
    SS12[30][40] = 4'hE;
    SS12[31][40] = 4'hE;
    SS12[32][40] = 4'h0;
    SS12[33][40] = 4'h0;
    SS12[34][40] = 4'h0;
    SS12[35][40] = 4'h0;
    SS12[36][40] = 4'h0;
    SS12[37][40] = 4'h0;
    SS12[38][40] = 4'h0;
    SS12[39][40] = 4'h0;
    SS12[40][40] = 4'h0;
    SS12[41][40] = 4'h0;
    SS12[42][40] = 4'h0;
    SS12[43][40] = 4'h0;
    SS12[44][40] = 4'h0;
    SS12[45][40] = 4'h0;
    SS12[46][40] = 4'h0;
    SS12[47][40] = 4'h0;
    SS12[0][41] = 4'h0;
    SS12[1][41] = 4'h0;
    SS12[2][41] = 4'h0;
    SS12[3][41] = 4'h0;
    SS12[4][41] = 4'h0;
    SS12[5][41] = 4'h0;
    SS12[6][41] = 4'h0;
    SS12[7][41] = 4'h0;
    SS12[8][41] = 4'h0;
    SS12[9][41] = 4'h0;
    SS12[10][41] = 4'h0;
    SS12[11][41] = 4'h0;
    SS12[12][41] = 4'hD;
    SS12[13][41] = 4'hD;
    SS12[14][41] = 4'hD;
    SS12[15][41] = 4'hD;
    SS12[16][41] = 4'hE;
    SS12[17][41] = 4'hE;
    SS12[18][41] = 4'hE;
    SS12[19][41] = 4'h0;
    SS12[20][41] = 4'h0;
    SS12[21][41] = 4'h0;
    SS12[22][41] = 4'h0;
    SS12[23][41] = 4'h0;
    SS12[24][41] = 4'h0;
    SS12[25][41] = 4'hC;
    SS12[26][41] = 4'hC;
    SS12[27][41] = 4'hC;
    SS12[28][41] = 4'hC;
    SS12[29][41] = 4'hE;
    SS12[30][41] = 4'hE;
    SS12[31][41] = 4'hE;
    SS12[32][41] = 4'h0;
    SS12[33][41] = 4'h0;
    SS12[34][41] = 4'h0;
    SS12[35][41] = 4'h0;
    SS12[36][41] = 4'h0;
    SS12[37][41] = 4'h0;
    SS12[38][41] = 4'h0;
    SS12[39][41] = 4'h0;
    SS12[40][41] = 4'h0;
    SS12[41][41] = 4'h0;
    SS12[42][41] = 4'h0;
    SS12[43][41] = 4'h0;
    SS12[44][41] = 4'h0;
    SS12[45][41] = 4'h0;
    SS12[46][41] = 4'h0;
    SS12[47][41] = 4'h0;
    SS12[0][42] = 4'h0;
    SS12[1][42] = 4'h0;
    SS12[2][42] = 4'h0;
    SS12[3][42] = 4'h0;
    SS12[4][42] = 4'h0;
    SS12[5][42] = 4'h0;
    SS12[6][42] = 4'h0;
    SS12[7][42] = 4'h0;
    SS12[8][42] = 4'h0;
    SS12[9][42] = 4'h0;
    SS12[10][42] = 4'h0;
    SS12[11][42] = 4'h0;
    SS12[12][42] = 4'h0;
    SS12[13][42] = 4'hD;
    SS12[14][42] = 4'hD;
    SS12[15][42] = 4'hD;
    SS12[16][42] = 4'hD;
    SS12[17][42] = 4'hE;
    SS12[18][42] = 4'h0;
    SS12[19][42] = 4'h0;
    SS12[20][42] = 4'h0;
    SS12[21][42] = 4'h0;
    SS12[22][42] = 4'h0;
    SS12[23][42] = 4'h0;
    SS12[24][42] = 4'h0;
    SS12[25][42] = 4'h0;
    SS12[26][42] = 4'hC;
    SS12[27][42] = 4'hC;
    SS12[28][42] = 4'hC;
    SS12[29][42] = 4'hC;
    SS12[30][42] = 4'hE;
    SS12[31][42] = 4'h0;
    SS12[32][42] = 4'h0;
    SS12[33][42] = 4'h0;
    SS12[34][42] = 4'h0;
    SS12[35][42] = 4'h0;
    SS12[36][42] = 4'h0;
    SS12[37][42] = 4'h0;
    SS12[38][42] = 4'h0;
    SS12[39][42] = 4'h0;
    SS12[40][42] = 4'h0;
    SS12[41][42] = 4'h0;
    SS12[42][42] = 4'h0;
    SS12[43][42] = 4'h0;
    SS12[44][42] = 4'h0;
    SS12[45][42] = 4'h0;
    SS12[46][42] = 4'h0;
    SS12[47][42] = 4'h0;
    SS12[0][43] = 4'h0;
    SS12[1][43] = 4'h0;
    SS12[2][43] = 4'h0;
    SS12[3][43] = 4'h0;
    SS12[4][43] = 4'h0;
    SS12[5][43] = 4'h0;
    SS12[6][43] = 4'h0;
    SS12[7][43] = 4'h0;
    SS12[8][43] = 4'h0;
    SS12[9][43] = 4'h0;
    SS12[10][43] = 4'h0;
    SS12[11][43] = 4'h0;
    SS12[12][43] = 4'h0;
    SS12[13][43] = 4'hD;
    SS12[14][43] = 4'hD;
    SS12[15][43] = 4'hD;
    SS12[16][43] = 4'hD;
    SS12[17][43] = 4'h0;
    SS12[18][43] = 4'h0;
    SS12[19][43] = 4'h0;
    SS12[20][43] = 4'h0;
    SS12[21][43] = 4'h0;
    SS12[22][43] = 4'h0;
    SS12[23][43] = 4'h0;
    SS12[24][43] = 4'h0;
    SS12[25][43] = 4'h0;
    SS12[26][43] = 4'hC;
    SS12[27][43] = 4'hC;
    SS12[28][43] = 4'hC;
    SS12[29][43] = 4'hC;
    SS12[30][43] = 4'hD;
    SS12[31][43] = 4'h0;
    SS12[32][43] = 4'h0;
    SS12[33][43] = 4'h0;
    SS12[34][43] = 4'h0;
    SS12[35][43] = 4'h0;
    SS12[36][43] = 4'h0;
    SS12[37][43] = 4'h0;
    SS12[38][43] = 4'h0;
    SS12[39][43] = 4'h0;
    SS12[40][43] = 4'h0;
    SS12[41][43] = 4'h0;
    SS12[42][43] = 4'h0;
    SS12[43][43] = 4'h0;
    SS12[44][43] = 4'h0;
    SS12[45][43] = 4'h0;
    SS12[46][43] = 4'h0;
    SS12[47][43] = 4'h0;
    SS12[0][44] = 4'h0;
    SS12[1][44] = 4'h0;
    SS12[2][44] = 4'h0;
    SS12[3][44] = 4'h0;
    SS12[4][44] = 4'h0;
    SS12[5][44] = 4'h0;
    SS12[6][44] = 4'h0;
    SS12[7][44] = 4'h0;
    SS12[8][44] = 4'h0;
    SS12[9][44] = 4'h0;
    SS12[10][44] = 4'h0;
    SS12[11][44] = 4'h0;
    SS12[12][44] = 4'hD;
    SS12[13][44] = 4'hD;
    SS12[14][44] = 4'hD;
    SS12[15][44] = 4'hD;
    SS12[16][44] = 4'h0;
    SS12[17][44] = 4'h0;
    SS12[18][44] = 4'h0;
    SS12[19][44] = 4'h0;
    SS12[20][44] = 4'h0;
    SS12[21][44] = 4'h0;
    SS12[22][44] = 4'h0;
    SS12[23][44] = 4'h0;
    SS12[24][44] = 4'h0;
    SS12[25][44] = 4'hC;
    SS12[26][44] = 4'hC;
    SS12[27][44] = 4'hC;
    SS12[28][44] = 4'hC;
    SS12[29][44] = 4'hD;
    SS12[30][44] = 4'hD;
    SS12[31][44] = 4'hD;
    SS12[32][44] = 4'h0;
    SS12[33][44] = 4'h0;
    SS12[34][44] = 4'h0;
    SS12[35][44] = 4'h0;
    SS12[36][44] = 4'h0;
    SS12[37][44] = 4'h0;
    SS12[38][44] = 4'h0;
    SS12[39][44] = 4'h0;
    SS12[40][44] = 4'h0;
    SS12[41][44] = 4'h0;
    SS12[42][44] = 4'h0;
    SS12[43][44] = 4'h0;
    SS12[44][44] = 4'h0;
    SS12[45][44] = 4'h0;
    SS12[46][44] = 4'h0;
    SS12[47][44] = 4'h0;
    SS12[0][45] = 4'h0;
    SS12[1][45] = 4'h0;
    SS12[2][45] = 4'h0;
    SS12[3][45] = 4'h0;
    SS12[4][45] = 4'h0;
    SS12[5][45] = 4'h0;
    SS12[6][45] = 4'h0;
    SS12[7][45] = 4'h0;
    SS12[8][45] = 4'h0;
    SS12[9][45] = 4'h0;
    SS12[10][45] = 4'h0;
    SS12[11][45] = 4'h0;
    SS12[12][45] = 4'hD;
    SS12[13][45] = 4'hD;
    SS12[14][45] = 4'hD;
    SS12[15][45] = 4'h0;
    SS12[16][45] = 4'h0;
    SS12[17][45] = 4'h0;
    SS12[18][45] = 4'h0;
    SS12[19][45] = 4'h0;
    SS12[20][45] = 4'h0;
    SS12[21][45] = 4'h0;
    SS12[22][45] = 4'h0;
    SS12[23][45] = 4'h0;
    SS12[24][45] = 4'hC;
    SS12[25][45] = 4'hC;
    SS12[26][45] = 4'hC;
    SS12[27][45] = 4'hC;
    SS12[28][45] = 4'hC;
    SS12[29][45] = 4'hD;
    SS12[30][45] = 4'hD;
    SS12[31][45] = 4'hD;
    SS12[32][45] = 4'h0;
    SS12[33][45] = 4'h0;
    SS12[34][45] = 4'h0;
    SS12[35][45] = 4'h0;
    SS12[36][45] = 4'h0;
    SS12[37][45] = 4'h0;
    SS12[38][45] = 4'h0;
    SS12[39][45] = 4'h0;
    SS12[40][45] = 4'h0;
    SS12[41][45] = 4'h0;
    SS12[42][45] = 4'h0;
    SS12[43][45] = 4'h0;
    SS12[44][45] = 4'h0;
    SS12[45][45] = 4'h0;
    SS12[46][45] = 4'h0;
    SS12[47][45] = 4'h0;
    SS12[0][46] = 4'h0;
    SS12[1][46] = 4'h0;
    SS12[2][46] = 4'h0;
    SS12[3][46] = 4'h0;
    SS12[4][46] = 4'h0;
    SS12[5][46] = 4'h0;
    SS12[6][46] = 4'h0;
    SS12[7][46] = 4'h0;
    SS12[8][46] = 4'h0;
    SS12[9][46] = 4'h0;
    SS12[10][46] = 4'h0;
    SS12[11][46] = 4'h0;
    SS12[12][46] = 4'h0;
    SS12[13][46] = 4'hD;
    SS12[14][46] = 4'h0;
    SS12[15][46] = 4'h0;
    SS12[16][46] = 4'h0;
    SS12[17][46] = 4'h0;
    SS12[18][46] = 4'h0;
    SS12[19][46] = 4'h0;
    SS12[20][46] = 4'h0;
    SS12[21][46] = 4'h0;
    SS12[22][46] = 4'h0;
    SS12[23][46] = 4'h0;
    SS12[24][46] = 4'h0;
    SS12[25][46] = 4'hC;
    SS12[26][46] = 4'hC;
    SS12[27][46] = 4'hC;
    SS12[28][46] = 4'hC;
    SS12[29][46] = 4'hC;
    SS12[30][46] = 4'hD;
    SS12[31][46] = 4'h0;
    SS12[32][46] = 4'h0;
    SS12[33][46] = 4'h0;
    SS12[34][46] = 4'h0;
    SS12[35][46] = 4'h0;
    SS12[36][46] = 4'h0;
    SS12[37][46] = 4'h0;
    SS12[38][46] = 4'h0;
    SS12[39][46] = 4'h0;
    SS12[40][46] = 4'h0;
    SS12[41][46] = 4'h0;
    SS12[42][46] = 4'h0;
    SS12[43][46] = 4'h0;
    SS12[44][46] = 4'h0;
    SS12[45][46] = 4'h0;
    SS12[46][46] = 4'h0;
    SS12[47][46] = 4'h0;
    SS12[0][47] = 4'h0;
    SS12[1][47] = 4'h0;
    SS12[2][47] = 4'h0;
    SS12[3][47] = 4'h0;
    SS12[4][47] = 4'h0;
    SS12[5][47] = 4'h0;
    SS12[6][47] = 4'h0;
    SS12[7][47] = 4'h0;
    SS12[8][47] = 4'h0;
    SS12[9][47] = 4'h0;
    SS12[10][47] = 4'h0;
    SS12[11][47] = 4'h0;
    SS12[12][47] = 4'h0;
    SS12[13][47] = 4'h0;
    SS12[14][47] = 4'h0;
    SS12[15][47] = 4'h0;
    SS12[16][47] = 4'h0;
    SS12[17][47] = 4'h0;
    SS12[18][47] = 4'h0;
    SS12[19][47] = 4'h0;
    SS12[20][47] = 4'h0;
    SS12[21][47] = 4'h0;
    SS12[22][47] = 4'h0;
    SS12[23][47] = 4'h0;
    SS12[24][47] = 4'h0;
    SS12[25][47] = 4'h0;
    SS12[26][47] = 4'hC;
    SS12[27][47] = 4'hC;
    SS12[28][47] = 4'hC;
    SS12[29][47] = 4'hC;
    SS12[30][47] = 4'hE;
    SS12[31][47] = 4'h0;
    SS12[32][47] = 4'h0;
    SS12[33][47] = 4'h0;
    SS12[34][47] = 4'h0;
    SS12[35][47] = 4'h0;
    SS12[36][47] = 4'h0;
    SS12[37][47] = 4'h0;
    SS12[38][47] = 4'h0;
    SS12[39][47] = 4'h0;
    SS12[40][47] = 4'h0;
    SS12[41][47] = 4'h0;
    SS12[42][47] = 4'h0;
    SS12[43][47] = 4'h0;
    SS12[44][47] = 4'h0;
    SS12[45][47] = 4'h0;
    SS12[46][47] = 4'h0;
    SS12[47][47] = 4'h0;
 
//SS 13
    SS13[0][0] = 4'h0;
    SS13[1][0] = 4'h0;
    SS13[2][0] = 4'h0;
    SS13[3][0] = 4'h0;
    SS13[4][0] = 4'h0;
    SS13[5][0] = 4'h0;
    SS13[6][0] = 4'h0;
    SS13[7][0] = 4'h0;
    SS13[8][0] = 4'h0;
    SS13[9][0] = 4'h0;
    SS13[10][0] = 4'h0;
    SS13[11][0] = 4'h0;
    SS13[12][0] = 4'h0;
    SS13[13][0] = 4'h0;
    SS13[14][0] = 4'h0;
    SS13[15][0] = 4'h0;
    SS13[16][0] = 4'h0;
    SS13[17][0] = 4'h0;
    SS13[18][0] = 4'h0;
    SS13[19][0] = 4'h0;
    SS13[20][0] = 4'h0;
    SS13[21][0] = 4'h0;
    SS13[22][0] = 4'h0;
    SS13[23][0] = 4'h0;
    SS13[24][0] = 4'h0;
    SS13[25][0] = 4'h0;
    SS13[26][0] = 4'h0;
    SS13[27][0] = 4'h0;
    SS13[28][0] = 4'h0;
    SS13[29][0] = 4'h0;
    SS13[30][0] = 4'h0;
    SS13[31][0] = 4'h0;
    SS13[32][0] = 4'h0;
    SS13[33][0] = 4'h0;
    SS13[34][0] = 4'h0;
    SS13[35][0] = 4'h0;
    SS13[36][0] = 4'h0;
    SS13[37][0] = 4'h0;
    SS13[38][0] = 4'h0;
    SS13[39][0] = 4'h0;
    SS13[40][0] = 4'h0;
    SS13[41][0] = 4'h0;
    SS13[42][0] = 4'h0;
    SS13[43][0] = 4'h0;
    SS13[44][0] = 4'h0;
    SS13[45][0] = 4'h0;
    SS13[46][0] = 4'h0;
    SS13[47][0] = 4'h0;
    SS13[0][1] = 4'h0;
    SS13[1][1] = 4'h0;
    SS13[2][1] = 4'h0;
    SS13[3][1] = 4'h0;
    SS13[4][1] = 4'h0;
    SS13[5][1] = 4'h0;
    SS13[6][1] = 4'h0;
    SS13[7][1] = 4'h0;
    SS13[8][1] = 4'h0;
    SS13[9][1] = 4'h0;
    SS13[10][1] = 4'h0;
    SS13[11][1] = 4'h0;
    SS13[12][1] = 4'h0;
    SS13[13][1] = 4'h0;
    SS13[14][1] = 4'h0;
    SS13[15][1] = 4'h0;
    SS13[16][1] = 4'hC;
    SS13[17][1] = 4'hC;
    SS13[18][1] = 4'h0;
    SS13[19][1] = 4'h0;
    SS13[20][1] = 4'h0;
    SS13[21][1] = 4'h0;
    SS13[22][1] = 4'h0;
    SS13[23][1] = 4'h0;
    SS13[24][1] = 4'h0;
    SS13[25][1] = 4'h0;
    SS13[26][1] = 4'h0;
    SS13[27][1] = 4'h0;
    SS13[28][1] = 4'h0;
    SS13[29][1] = 4'h0;
    SS13[30][1] = 4'h0;
    SS13[31][1] = 4'h0;
    SS13[32][1] = 4'h0;
    SS13[33][1] = 4'h0;
    SS13[34][1] = 4'h0;
    SS13[35][1] = 4'h0;
    SS13[36][1] = 4'h0;
    SS13[37][1] = 4'h0;
    SS13[38][1] = 4'h0;
    SS13[39][1] = 4'h0;
    SS13[40][1] = 4'h0;
    SS13[41][1] = 4'h0;
    SS13[42][1] = 4'h0;
    SS13[43][1] = 4'h0;
    SS13[44][1] = 4'h0;
    SS13[45][1] = 4'h0;
    SS13[46][1] = 4'h0;
    SS13[47][1] = 4'h0;
    SS13[0][2] = 4'h0;
    SS13[1][2] = 4'h0;
    SS13[2][2] = 4'h0;
    SS13[3][2] = 4'h0;
    SS13[4][2] = 4'h0;
    SS13[5][2] = 4'h0;
    SS13[6][2] = 4'h0;
    SS13[7][2] = 4'h0;
    SS13[8][2] = 4'h0;
    SS13[9][2] = 4'h0;
    SS13[10][2] = 4'h0;
    SS13[11][2] = 4'h0;
    SS13[12][2] = 4'h0;
    SS13[13][2] = 4'h0;
    SS13[14][2] = 4'hC;
    SS13[15][2] = 4'hC;
    SS13[16][2] = 4'hC;
    SS13[17][2] = 4'hC;
    SS13[18][2] = 4'h0;
    SS13[19][2] = 4'h0;
    SS13[20][2] = 4'h0;
    SS13[21][2] = 4'h0;
    SS13[22][2] = 4'h0;
    SS13[23][2] = 4'h0;
    SS13[24][2] = 4'h0;
    SS13[25][2] = 4'h0;
    SS13[26][2] = 4'h0;
    SS13[27][2] = 4'h0;
    SS13[28][2] = 4'h0;
    SS13[29][2] = 4'h0;
    SS13[30][2] = 4'h0;
    SS13[31][2] = 4'h0;
    SS13[32][2] = 4'h0;
    SS13[33][2] = 4'h0;
    SS13[34][2] = 4'h0;
    SS13[35][2] = 4'h0;
    SS13[36][2] = 4'h0;
    SS13[37][2] = 4'h0;
    SS13[38][2] = 4'h0;
    SS13[39][2] = 4'h0;
    SS13[40][2] = 4'h0;
    SS13[41][2] = 4'h0;
    SS13[42][2] = 4'h0;
    SS13[43][2] = 4'h0;
    SS13[44][2] = 4'h0;
    SS13[45][2] = 4'h0;
    SS13[46][2] = 4'h0;
    SS13[47][2] = 4'h0;
    SS13[0][3] = 4'h0;
    SS13[1][3] = 4'h0;
    SS13[2][3] = 4'h0;
    SS13[3][3] = 4'h0;
    SS13[4][3] = 4'h0;
    SS13[5][3] = 4'h0;
    SS13[6][3] = 4'h0;
    SS13[7][3] = 4'h0;
    SS13[8][3] = 4'h0;
    SS13[9][3] = 4'h0;
    SS13[10][3] = 4'h0;
    SS13[11][3] = 4'h0;
    SS13[12][3] = 4'hC;
    SS13[13][3] = 4'hC;
    SS13[14][3] = 4'hC;
    SS13[15][3] = 4'hC;
    SS13[16][3] = 4'hC;
    SS13[17][3] = 4'hC;
    SS13[18][3] = 4'hC;
    SS13[19][3] = 4'h0;
    SS13[20][3] = 4'h0;
    SS13[21][3] = 4'h0;
    SS13[22][3] = 4'h0;
    SS13[23][3] = 4'h0;
    SS13[24][3] = 4'h0;
    SS13[25][3] = 4'h0;
    SS13[26][3] = 4'h0;
    SS13[27][3] = 4'h0;
    SS13[28][3] = 4'h0;
    SS13[29][3] = 4'h0;
    SS13[30][3] = 4'h0;
    SS13[31][3] = 4'h0;
    SS13[32][3] = 4'h0;
    SS13[33][3] = 4'h0;
    SS13[34][3] = 4'h0;
    SS13[35][3] = 4'h0;
    SS13[36][3] = 4'h0;
    SS13[37][3] = 4'h0;
    SS13[38][3] = 4'h0;
    SS13[39][3] = 4'h0;
    SS13[40][3] = 4'h0;
    SS13[41][3] = 4'h0;
    SS13[42][3] = 4'h0;
    SS13[43][3] = 4'h0;
    SS13[44][3] = 4'h0;
    SS13[45][3] = 4'h0;
    SS13[46][3] = 4'h0;
    SS13[47][3] = 4'h0;
    SS13[0][4] = 4'h0;
    SS13[1][4] = 4'h0;
    SS13[2][4] = 4'h0;
    SS13[3][4] = 4'h0;
    SS13[4][4] = 4'h0;
    SS13[5][4] = 4'h0;
    SS13[6][4] = 4'h0;
    SS13[7][4] = 4'h0;
    SS13[8][4] = 4'h0;
    SS13[9][4] = 4'h0;
    SS13[10][4] = 4'h0;
    SS13[11][4] = 4'h0;
    SS13[12][4] = 4'h0;
    SS13[13][4] = 4'hC;
    SS13[14][4] = 4'hC;
    SS13[15][4] = 4'hC;
    SS13[16][4] = 4'hC;
    SS13[17][4] = 4'hC;
    SS13[18][4] = 4'hC;
    SS13[19][4] = 4'h0;
    SS13[20][4] = 4'h0;
    SS13[21][4] = 4'h0;
    SS13[22][4] = 4'h0;
    SS13[23][4] = 4'h0;
    SS13[24][4] = 4'h0;
    SS13[25][4] = 4'h0;
    SS13[26][4] = 4'h0;
    SS13[27][4] = 4'h0;
    SS13[28][4] = 4'h0;
    SS13[29][4] = 4'h0;
    SS13[30][4] = 4'h0;
    SS13[31][4] = 4'h0;
    SS13[32][4] = 4'h0;
    SS13[33][4] = 4'h0;
    SS13[34][4] = 4'h0;
    SS13[35][4] = 4'h0;
    SS13[36][4] = 4'h0;
    SS13[37][4] = 4'h0;
    SS13[38][4] = 4'h0;
    SS13[39][4] = 4'h0;
    SS13[40][4] = 4'h0;
    SS13[41][4] = 4'h0;
    SS13[42][4] = 4'h0;
    SS13[43][4] = 4'h0;
    SS13[44][4] = 4'h0;
    SS13[45][4] = 4'h0;
    SS13[46][4] = 4'h0;
    SS13[47][4] = 4'h0;
    SS13[0][5] = 4'h0;
    SS13[1][5] = 4'h0;
    SS13[2][5] = 4'h0;
    SS13[3][5] = 4'h0;
    SS13[4][5] = 4'h0;
    SS13[5][5] = 4'h0;
    SS13[6][5] = 4'h0;
    SS13[7][5] = 4'h0;
    SS13[8][5] = 4'h0;
    SS13[9][5] = 4'h0;
    SS13[10][5] = 4'h0;
    SS13[11][5] = 4'h0;
    SS13[12][5] = 4'h0;
    SS13[13][5] = 4'hC;
    SS13[14][5] = 4'hC;
    SS13[15][5] = 4'hC;
    SS13[16][5] = 4'hC;
    SS13[17][5] = 4'hC;
    SS13[18][5] = 4'hC;
    SS13[19][5] = 4'hC;
    SS13[20][5] = 4'h0;
    SS13[21][5] = 4'h0;
    SS13[22][5] = 4'hD;
    SS13[23][5] = 4'h0;
    SS13[24][5] = 4'h0;
    SS13[25][5] = 4'h0;
    SS13[26][5] = 4'h0;
    SS13[27][5] = 4'h0;
    SS13[28][5] = 4'h0;
    SS13[29][5] = 4'h0;
    SS13[30][5] = 4'h0;
    SS13[31][5] = 4'h0;
    SS13[32][5] = 4'h0;
    SS13[33][5] = 4'h0;
    SS13[34][5] = 4'h0;
    SS13[35][5] = 4'h0;
    SS13[36][5] = 4'h0;
    SS13[37][5] = 4'h0;
    SS13[38][5] = 4'h0;
    SS13[39][5] = 4'h0;
    SS13[40][5] = 4'h0;
    SS13[41][5] = 4'h0;
    SS13[42][5] = 4'h0;
    SS13[43][5] = 4'h0;
    SS13[44][5] = 4'h0;
    SS13[45][5] = 4'h0;
    SS13[46][5] = 4'h0;
    SS13[47][5] = 4'h0;
    SS13[0][6] = 4'h0;
    SS13[1][6] = 4'h0;
    SS13[2][6] = 4'h0;
    SS13[3][6] = 4'h0;
    SS13[4][6] = 4'h0;
    SS13[5][6] = 4'h0;
    SS13[6][6] = 4'h0;
    SS13[7][6] = 4'h0;
    SS13[8][6] = 4'h0;
    SS13[9][6] = 4'h0;
    SS13[10][6] = 4'h0;
    SS13[11][6] = 4'h0;
    SS13[12][6] = 4'h0;
    SS13[13][6] = 4'h0;
    SS13[14][6] = 4'hC;
    SS13[15][6] = 4'hC;
    SS13[16][6] = 4'hC;
    SS13[17][6] = 4'hC;
    SS13[18][6] = 4'hC;
    SS13[19][6] = 4'hC;
    SS13[20][6] = 4'hD;
    SS13[21][6] = 4'hD;
    SS13[22][6] = 4'hD;
    SS13[23][6] = 4'h0;
    SS13[24][6] = 4'h0;
    SS13[25][6] = 4'h0;
    SS13[26][6] = 4'h0;
    SS13[27][6] = 4'h0;
    SS13[28][6] = 4'h0;
    SS13[29][6] = 4'h0;
    SS13[30][6] = 4'h0;
    SS13[31][6] = 4'h0;
    SS13[32][6] = 4'h0;
    SS13[33][6] = 4'h0;
    SS13[34][6] = 4'h0;
    SS13[35][6] = 4'h0;
    SS13[36][6] = 4'h0;
    SS13[37][6] = 4'h0;
    SS13[38][6] = 4'h0;
    SS13[39][6] = 4'h0;
    SS13[40][6] = 4'h0;
    SS13[41][6] = 4'h0;
    SS13[42][6] = 4'h0;
    SS13[43][6] = 4'h0;
    SS13[44][6] = 4'h0;
    SS13[45][6] = 4'h0;
    SS13[46][6] = 4'h0;
    SS13[47][6] = 4'h0;
    SS13[0][7] = 4'h0;
    SS13[1][7] = 4'h0;
    SS13[2][7] = 4'h0;
    SS13[3][7] = 4'h0;
    SS13[4][7] = 4'h0;
    SS13[5][7] = 4'h0;
    SS13[6][7] = 4'h0;
    SS13[7][7] = 4'h0;
    SS13[8][7] = 4'h0;
    SS13[9][7] = 4'h0;
    SS13[10][7] = 4'h0;
    SS13[11][7] = 4'h0;
    SS13[12][7] = 4'h0;
    SS13[13][7] = 4'h0;
    SS13[14][7] = 4'hC;
    SS13[15][7] = 4'hC;
    SS13[16][7] = 4'hC;
    SS13[17][7] = 4'hC;
    SS13[18][7] = 4'hC;
    SS13[19][7] = 4'hC;
    SS13[20][7] = 4'hD;
    SS13[21][7] = 4'hD;
    SS13[22][7] = 4'hD;
    SS13[23][7] = 4'hD;
    SS13[24][7] = 4'h0;
    SS13[25][7] = 4'h0;
    SS13[26][7] = 4'h0;
    SS13[27][7] = 4'h0;
    SS13[28][7] = 4'h0;
    SS13[29][7] = 4'h0;
    SS13[30][7] = 4'h0;
    SS13[31][7] = 4'h0;
    SS13[32][7] = 4'h0;
    SS13[33][7] = 4'h0;
    SS13[34][7] = 4'h0;
    SS13[35][7] = 4'h0;
    SS13[36][7] = 4'h0;
    SS13[37][7] = 4'h0;
    SS13[38][7] = 4'h0;
    SS13[39][7] = 4'h0;
    SS13[40][7] = 4'h0;
    SS13[41][7] = 4'h0;
    SS13[42][7] = 4'h0;
    SS13[43][7] = 4'h0;
    SS13[44][7] = 4'h0;
    SS13[45][7] = 4'h0;
    SS13[46][7] = 4'h0;
    SS13[47][7] = 4'h0;
    SS13[0][8] = 4'h0;
    SS13[1][8] = 4'h0;
    SS13[2][8] = 4'h0;
    SS13[3][8] = 4'h0;
    SS13[4][8] = 4'h0;
    SS13[5][8] = 4'h0;
    SS13[6][8] = 4'h0;
    SS13[7][8] = 4'h0;
    SS13[8][8] = 4'h0;
    SS13[9][8] = 4'h0;
    SS13[10][8] = 4'h0;
    SS13[11][8] = 4'h0;
    SS13[12][8] = 4'h0;
    SS13[13][8] = 4'h0;
    SS13[14][8] = 4'hC;
    SS13[15][8] = 4'hC;
    SS13[16][8] = 4'hC;
    SS13[17][8] = 4'hC;
    SS13[18][8] = 4'hC;
    SS13[19][8] = 4'hC;
    SS13[20][8] = 4'hC;
    SS13[21][8] = 4'hD;
    SS13[22][8] = 4'hD;
    SS13[23][8] = 4'hD;
    SS13[24][8] = 4'h0;
    SS13[25][8] = 4'h0;
    SS13[26][8] = 4'h0;
    SS13[27][8] = 4'h0;
    SS13[28][8] = 4'h0;
    SS13[29][8] = 4'h0;
    SS13[30][8] = 4'h0;
    SS13[31][8] = 4'h0;
    SS13[32][8] = 4'h0;
    SS13[33][8] = 4'h0;
    SS13[34][8] = 4'h0;
    SS13[35][8] = 4'h0;
    SS13[36][8] = 4'h0;
    SS13[37][8] = 4'h0;
    SS13[38][8] = 4'h0;
    SS13[39][8] = 4'h0;
    SS13[40][8] = 4'h0;
    SS13[41][8] = 4'h0;
    SS13[42][8] = 4'h0;
    SS13[43][8] = 4'h0;
    SS13[44][8] = 4'h0;
    SS13[45][8] = 4'h0;
    SS13[46][8] = 4'h0;
    SS13[47][8] = 4'h0;
    SS13[0][9] = 4'h0;
    SS13[1][9] = 4'h0;
    SS13[2][9] = 4'h0;
    SS13[3][9] = 4'h0;
    SS13[4][9] = 4'h0;
    SS13[5][9] = 4'h0;
    SS13[6][9] = 4'h0;
    SS13[7][9] = 4'h0;
    SS13[8][9] = 4'h0;
    SS13[9][9] = 4'h0;
    SS13[10][9] = 4'h0;
    SS13[11][9] = 4'h0;
    SS13[12][9] = 4'hF;
    SS13[13][9] = 4'hD;
    SS13[14][9] = 4'hD;
    SS13[15][9] = 4'hC;
    SS13[16][9] = 4'hC;
    SS13[17][9] = 4'hC;
    SS13[18][9] = 4'hC;
    SS13[19][9] = 4'hC;
    SS13[20][9] = 4'hC;
    SS13[21][9] = 4'hD;
    SS13[22][9] = 4'hD;
    SS13[23][9] = 4'hD;
    SS13[24][9] = 4'h0;
    SS13[25][9] = 4'h0;
    SS13[26][9] = 4'h0;
    SS13[27][9] = 4'h0;
    SS13[28][9] = 4'h0;
    SS13[29][9] = 4'h0;
    SS13[30][9] = 4'h0;
    SS13[31][9] = 4'h0;
    SS13[32][9] = 4'h0;
    SS13[33][9] = 4'h0;
    SS13[34][9] = 4'h0;
    SS13[35][9] = 4'h0;
    SS13[36][9] = 4'h0;
    SS13[37][9] = 4'h0;
    SS13[38][9] = 4'h0;
    SS13[39][9] = 4'h0;
    SS13[40][9] = 4'h0;
    SS13[41][9] = 4'h0;
    SS13[42][9] = 4'h0;
    SS13[43][9] = 4'h0;
    SS13[44][9] = 4'h0;
    SS13[45][9] = 4'h0;
    SS13[46][9] = 4'h0;
    SS13[47][9] = 4'h0;
    SS13[0][10] = 4'h0;
    SS13[1][10] = 4'h0;
    SS13[2][10] = 4'h0;
    SS13[3][10] = 4'h0;
    SS13[4][10] = 4'h0;
    SS13[5][10] = 4'h0;
    SS13[6][10] = 4'h0;
    SS13[7][10] = 4'h0;
    SS13[8][10] = 4'h0;
    SS13[9][10] = 4'h0;
    SS13[10][10] = 4'h0;
    SS13[11][10] = 4'h0;
    SS13[12][10] = 4'hD;
    SS13[13][10] = 4'hD;
    SS13[14][10] = 4'hD;
    SS13[15][10] = 4'hC;
    SS13[16][10] = 4'hC;
    SS13[17][10] = 4'hC;
    SS13[18][10] = 4'hC;
    SS13[19][10] = 4'hC;
    SS13[20][10] = 4'hC;
    SS13[21][10] = 4'hC;
    SS13[22][10] = 4'hD;
    SS13[23][10] = 4'hD;
    SS13[24][10] = 4'hD;
    SS13[25][10] = 4'h0;
    SS13[26][10] = 4'h0;
    SS13[27][10] = 4'h0;
    SS13[28][10] = 4'h0;
    SS13[29][10] = 4'h0;
    SS13[30][10] = 4'h0;
    SS13[31][10] = 4'h0;
    SS13[32][10] = 4'h0;
    SS13[33][10] = 4'h0;
    SS13[34][10] = 4'h0;
    SS13[35][10] = 4'h0;
    SS13[36][10] = 4'h0;
    SS13[37][10] = 4'h0;
    SS13[38][10] = 4'h0;
    SS13[39][10] = 4'h0;
    SS13[40][10] = 4'h0;
    SS13[41][10] = 4'h0;
    SS13[42][10] = 4'h0;
    SS13[43][10] = 4'h0;
    SS13[44][10] = 4'h0;
    SS13[45][10] = 4'h0;
    SS13[46][10] = 4'h0;
    SS13[47][10] = 4'h0;
    SS13[0][11] = 4'h0;
    SS13[1][11] = 4'h0;
    SS13[2][11] = 4'h0;
    SS13[3][11] = 4'h0;
    SS13[4][11] = 4'h0;
    SS13[5][11] = 4'h0;
    SS13[6][11] = 4'h0;
    SS13[7][11] = 4'h0;
    SS13[8][11] = 4'h0;
    SS13[9][11] = 4'h0;
    SS13[10][11] = 4'h0;
    SS13[11][11] = 4'h0;
    SS13[12][11] = 4'hD;
    SS13[13][11] = 4'hD;
    SS13[14][11] = 4'hD;
    SS13[15][11] = 4'hD;
    SS13[16][11] = 4'hC;
    SS13[17][11] = 4'hC;
    SS13[18][11] = 4'hC;
    SS13[19][11] = 4'hC;
    SS13[20][11] = 4'hC;
    SS13[21][11] = 4'hC;
    SS13[22][11] = 4'hD;
    SS13[23][11] = 4'hD;
    SS13[24][11] = 4'hD;
    SS13[25][11] = 4'h0;
    SS13[26][11] = 4'h0;
    SS13[27][11] = 4'h0;
    SS13[28][11] = 4'h0;
    SS13[29][11] = 4'h0;
    SS13[30][11] = 4'h0;
    SS13[31][11] = 4'h0;
    SS13[32][11] = 4'h0;
    SS13[33][11] = 4'h0;
    SS13[34][11] = 4'h0;
    SS13[35][11] = 4'h0;
    SS13[36][11] = 4'h0;
    SS13[37][11] = 4'h0;
    SS13[38][11] = 4'h0;
    SS13[39][11] = 4'h0;
    SS13[40][11] = 4'h0;
    SS13[41][11] = 4'h0;
    SS13[42][11] = 4'h0;
    SS13[43][11] = 4'h0;
    SS13[44][11] = 4'h0;
    SS13[45][11] = 4'h0;
    SS13[46][11] = 4'h0;
    SS13[47][11] = 4'h0;
    SS13[0][12] = 4'h0;
    SS13[1][12] = 4'h0;
    SS13[2][12] = 4'h0;
    SS13[3][12] = 4'h0;
    SS13[4][12] = 4'h0;
    SS13[5][12] = 4'h0;
    SS13[6][12] = 4'h0;
    SS13[7][12] = 4'h0;
    SS13[8][12] = 4'h0;
    SS13[9][12] = 4'h0;
    SS13[10][12] = 4'h0;
    SS13[11][12] = 4'h0;
    SS13[12][12] = 4'h0;
    SS13[13][12] = 4'hD;
    SS13[14][12] = 4'hD;
    SS13[15][12] = 4'hD;
    SS13[16][12] = 4'hC;
    SS13[17][12] = 4'hC;
    SS13[18][12] = 4'hC;
    SS13[19][12] = 4'hC;
    SS13[20][12] = 4'hC;
    SS13[21][12] = 4'hC;
    SS13[22][12] = 4'hD;
    SS13[23][12] = 4'hD;
    SS13[24][12] = 4'hD;
    SS13[25][12] = 4'hD;
    SS13[26][12] = 4'h0;
    SS13[27][12] = 4'h0;
    SS13[28][12] = 4'h0;
    SS13[29][12] = 4'h0;
    SS13[30][12] = 4'h0;
    SS13[31][12] = 4'h0;
    SS13[32][12] = 4'h0;
    SS13[33][12] = 4'h0;
    SS13[34][12] = 4'h0;
    SS13[35][12] = 4'h0;
    SS13[36][12] = 4'h0;
    SS13[37][12] = 4'h0;
    SS13[38][12] = 4'h0;
    SS13[39][12] = 4'h0;
    SS13[40][12] = 4'h0;
    SS13[41][12] = 4'h0;
    SS13[42][12] = 4'h0;
    SS13[43][12] = 4'h0;
    SS13[44][12] = 4'h0;
    SS13[45][12] = 4'h0;
    SS13[46][12] = 4'h0;
    SS13[47][12] = 4'h0;
    SS13[0][13] = 4'h0;
    SS13[1][13] = 4'h0;
    SS13[2][13] = 4'h0;
    SS13[3][13] = 4'h0;
    SS13[4][13] = 4'h0;
    SS13[5][13] = 4'h0;
    SS13[6][13] = 4'h0;
    SS13[7][13] = 4'h0;
    SS13[8][13] = 4'h0;
    SS13[9][13] = 4'h0;
    SS13[10][13] = 4'h0;
    SS13[11][13] = 4'h0;
    SS13[12][13] = 4'h0;
    SS13[13][13] = 4'hD;
    SS13[14][13] = 4'hD;
    SS13[15][13] = 4'hD;
    SS13[16][13] = 4'hC;
    SS13[17][13] = 4'hC;
    SS13[18][13] = 4'hC;
    SS13[19][13] = 4'hC;
    SS13[20][13] = 4'hC;
    SS13[21][13] = 4'hC;
    SS13[22][13] = 4'hC;
    SS13[23][13] = 4'hD;
    SS13[24][13] = 4'hD;
    SS13[25][13] = 4'hD;
    SS13[26][13] = 4'h0;
    SS13[27][13] = 4'h0;
    SS13[28][13] = 4'h0;
    SS13[29][13] = 4'h0;
    SS13[30][13] = 4'h0;
    SS13[31][13] = 4'h0;
    SS13[32][13] = 4'h0;
    SS13[33][13] = 4'h0;
    SS13[34][13] = 4'h0;
    SS13[35][13] = 4'h0;
    SS13[36][13] = 4'h0;
    SS13[37][13] = 4'h0;
    SS13[38][13] = 4'h0;
    SS13[39][13] = 4'h0;
    SS13[40][13] = 4'h0;
    SS13[41][13] = 4'h0;
    SS13[42][13] = 4'h0;
    SS13[43][13] = 4'h0;
    SS13[44][13] = 4'h0;
    SS13[45][13] = 4'h0;
    SS13[46][13] = 4'h0;
    SS13[47][13] = 4'h0;
    SS13[0][14] = 4'h0;
    SS13[1][14] = 4'h0;
    SS13[2][14] = 4'h0;
    SS13[3][14] = 4'h0;
    SS13[4][14] = 4'h0;
    SS13[5][14] = 4'h0;
    SS13[6][14] = 4'h0;
    SS13[7][14] = 4'h0;
    SS13[8][14] = 4'h0;
    SS13[9][14] = 4'h0;
    SS13[10][14] = 4'h0;
    SS13[11][14] = 4'h0;
    SS13[12][14] = 4'h0;
    SS13[13][14] = 4'h0;
    SS13[14][14] = 4'hD;
    SS13[15][14] = 4'hD;
    SS13[16][14] = 4'hD;
    SS13[17][14] = 4'hC;
    SS13[18][14] = 4'hC;
    SS13[19][14] = 4'hC;
    SS13[20][14] = 4'hC;
    SS13[21][14] = 4'hC;
    SS13[22][14] = 4'hC;
    SS13[23][14] = 4'hD;
    SS13[24][14] = 4'hC;
    SS13[25][14] = 4'hC;
    SS13[26][14] = 4'hE;
    SS13[27][14] = 4'h0;
    SS13[28][14] = 4'h0;
    SS13[29][14] = 4'h0;
    SS13[30][14] = 4'h0;
    SS13[31][14] = 4'h3;
    SS13[32][14] = 4'h3;
    SS13[33][14] = 4'h0;
    SS13[34][14] = 4'h0;
    SS13[35][14] = 4'h0;
    SS13[36][14] = 4'h0;
    SS13[37][14] = 4'h0;
    SS13[38][14] = 4'h0;
    SS13[39][14] = 4'h0;
    SS13[40][14] = 4'h0;
    SS13[41][14] = 4'h0;
    SS13[42][14] = 4'h0;
    SS13[43][14] = 4'h0;
    SS13[44][14] = 4'h0;
    SS13[45][14] = 4'h0;
    SS13[46][14] = 4'h0;
    SS13[47][14] = 4'h0;
    SS13[0][15] = 4'h0;
    SS13[1][15] = 4'h0;
    SS13[2][15] = 4'h0;
    SS13[3][15] = 4'h0;
    SS13[4][15] = 4'h0;
    SS13[5][15] = 4'h0;
    SS13[6][15] = 4'h0;
    SS13[7][15] = 4'h0;
    SS13[8][15] = 4'h0;
    SS13[9][15] = 4'h0;
    SS13[10][15] = 4'h0;
    SS13[11][15] = 4'h0;
    SS13[12][15] = 4'h0;
    SS13[13][15] = 4'h0;
    SS13[14][15] = 4'hD;
    SS13[15][15] = 4'hD;
    SS13[16][15] = 4'hD;
    SS13[17][15] = 4'hC;
    SS13[18][15] = 4'hC;
    SS13[19][15] = 4'hC;
    SS13[20][15] = 4'hC;
    SS13[21][15] = 4'hC;
    SS13[22][15] = 4'hC;
    SS13[23][15] = 4'hC;
    SS13[24][15] = 4'hC;
    SS13[25][15] = 4'hC;
    SS13[26][15] = 4'hC;
    SS13[27][15] = 4'h0;
    SS13[28][15] = 4'h0;
    SS13[29][15] = 4'hD;
    SS13[30][15] = 4'h3;
    SS13[31][15] = 4'h3;
    SS13[32][15] = 4'h3;
    SS13[33][15] = 4'h0;
    SS13[34][15] = 4'h0;
    SS13[35][15] = 4'h0;
    SS13[36][15] = 4'h0;
    SS13[37][15] = 4'h0;
    SS13[38][15] = 4'h0;
    SS13[39][15] = 4'h0;
    SS13[40][15] = 4'h0;
    SS13[41][15] = 4'h0;
    SS13[42][15] = 4'h0;
    SS13[43][15] = 4'h0;
    SS13[44][15] = 4'h0;
    SS13[45][15] = 4'h0;
    SS13[46][15] = 4'h0;
    SS13[47][15] = 4'h0;
    SS13[0][16] = 4'h0;
    SS13[1][16] = 4'h0;
    SS13[2][16] = 4'h0;
    SS13[3][16] = 4'h0;
    SS13[4][16] = 4'h0;
    SS13[5][16] = 4'h0;
    SS13[6][16] = 4'h0;
    SS13[7][16] = 4'h0;
    SS13[8][16] = 4'h0;
    SS13[9][16] = 4'h0;
    SS13[10][16] = 4'h0;
    SS13[11][16] = 4'h0;
    SS13[12][16] = 4'h0;
    SS13[13][16] = 4'h0;
    SS13[14][16] = 4'hD;
    SS13[15][16] = 4'hD;
    SS13[16][16] = 4'hD;
    SS13[17][16] = 4'hD;
    SS13[18][16] = 4'hC;
    SS13[19][16] = 4'hC;
    SS13[20][16] = 4'hC;
    SS13[21][16] = 4'hC;
    SS13[22][16] = 4'hC;
    SS13[23][16] = 4'hC;
    SS13[24][16] = 4'hC;
    SS13[25][16] = 4'hC;
    SS13[26][16] = 4'hC;
    SS13[27][16] = 4'hD;
    SS13[28][16] = 4'hD;
    SS13[29][16] = 4'hD;
    SS13[30][16] = 4'hD;
    SS13[31][16] = 4'h3;
    SS13[32][16] = 4'h3;
    SS13[33][16] = 4'h3;
    SS13[34][16] = 4'h0;
    SS13[35][16] = 4'h0;
    SS13[36][16] = 4'h0;
    SS13[37][16] = 4'h0;
    SS13[38][16] = 4'h0;
    SS13[39][16] = 4'h0;
    SS13[40][16] = 4'h0;
    SS13[41][16] = 4'h0;
    SS13[42][16] = 4'h0;
    SS13[43][16] = 4'h0;
    SS13[44][16] = 4'h0;
    SS13[45][16] = 4'h0;
    SS13[46][16] = 4'h0;
    SS13[47][16] = 4'h0;
    SS13[0][17] = 4'h0;
    SS13[1][17] = 4'h0;
    SS13[2][17] = 4'h0;
    SS13[3][17] = 4'h0;
    SS13[4][17] = 4'h0;
    SS13[5][17] = 4'h0;
    SS13[6][17] = 4'h0;
    SS13[7][17] = 4'h0;
    SS13[8][17] = 4'h0;
    SS13[9][17] = 4'h0;
    SS13[10][17] = 4'h0;
    SS13[11][17] = 4'h0;
    SS13[12][17] = 4'h0;
    SS13[13][17] = 4'h0;
    SS13[14][17] = 4'h0;
    SS13[15][17] = 4'hD;
    SS13[16][17] = 4'hC;
    SS13[17][17] = 4'hC;
    SS13[18][17] = 4'hC;
    SS13[19][17] = 4'hC;
    SS13[20][17] = 4'hC;
    SS13[21][17] = 4'hC;
    SS13[22][17] = 4'hC;
    SS13[23][17] = 4'hC;
    SS13[24][17] = 4'hA;
    SS13[25][17] = 4'hD;
    SS13[26][17] = 4'hD;
    SS13[27][17] = 4'hD;
    SS13[28][17] = 4'hD;
    SS13[29][17] = 4'hD;
    SS13[30][17] = 4'hD;
    SS13[31][17] = 4'h3;
    SS13[32][17] = 4'hD;
    SS13[33][17] = 4'hD;
    SS13[34][17] = 4'h0;
    SS13[35][17] = 4'h0;
    SS13[36][17] = 4'h0;
    SS13[37][17] = 4'h0;
    SS13[38][17] = 4'h0;
    SS13[39][17] = 4'h0;
    SS13[40][17] = 4'h3;
    SS13[41][17] = 4'h0;
    SS13[42][17] = 4'h0;
    SS13[43][17] = 4'h0;
    SS13[44][17] = 4'h0;
    SS13[45][17] = 4'h0;
    SS13[46][17] = 4'h0;
    SS13[47][17] = 4'h0;
    SS13[0][18] = 4'h0;
    SS13[1][18] = 4'h0;
    SS13[2][18] = 4'h0;
    SS13[3][18] = 4'h0;
    SS13[4][18] = 4'h0;
    SS13[5][18] = 4'h0;
    SS13[6][18] = 4'h0;
    SS13[7][18] = 4'h0;
    SS13[8][18] = 4'h0;
    SS13[9][18] = 4'h0;
    SS13[10][18] = 4'h0;
    SS13[11][18] = 4'h0;
    SS13[12][18] = 4'h0;
    SS13[13][18] = 4'h0;
    SS13[14][18] = 4'h0;
    SS13[15][18] = 4'hC;
    SS13[16][18] = 4'hC;
    SS13[17][18] = 4'hC;
    SS13[18][18] = 4'hC;
    SS13[19][18] = 4'hC;
    SS13[20][18] = 4'hC;
    SS13[21][18] = 4'hC;
    SS13[22][18] = 4'hA;
    SS13[23][18] = 4'hA;
    SS13[24][18] = 4'hA;
    SS13[25][18] = 4'hD;
    SS13[26][18] = 4'hD;
    SS13[27][18] = 4'hD;
    SS13[28][18] = 4'hD;
    SS13[29][18] = 4'hD;
    SS13[30][18] = 4'hD;
    SS13[31][18] = 4'hD;
    SS13[32][18] = 4'hD;
    SS13[33][18] = 4'hD;
    SS13[34][18] = 4'hD;
    SS13[35][18] = 4'h0;
    SS13[36][18] = 4'h0;
    SS13[37][18] = 4'hD;
    SS13[38][18] = 4'h3;
    SS13[39][18] = 4'h3;
    SS13[40][18] = 4'h3;
    SS13[41][18] = 4'h0;
    SS13[42][18] = 4'h0;
    SS13[43][18] = 4'h0;
    SS13[44][18] = 4'h0;
    SS13[45][18] = 4'h0;
    SS13[46][18] = 4'h0;
    SS13[47][18] = 4'h0;
    SS13[0][19] = 4'h0;
    SS13[1][19] = 4'h0;
    SS13[2][19] = 4'h0;
    SS13[3][19] = 4'h0;
    SS13[4][19] = 4'h0;
    SS13[5][19] = 4'h0;
    SS13[6][19] = 4'h0;
    SS13[7][19] = 4'h0;
    SS13[8][19] = 4'h0;
    SS13[9][19] = 4'h0;
    SS13[10][19] = 4'h0;
    SS13[11][19] = 4'h0;
    SS13[12][19] = 4'h0;
    SS13[13][19] = 4'h0;
    SS13[14][19] = 4'h0;
    SS13[15][19] = 4'h0;
    SS13[16][19] = 4'hC;
    SS13[17][19] = 4'hC;
    SS13[18][19] = 4'hC;
    SS13[19][19] = 4'hA;
    SS13[20][19] = 4'hA;
    SS13[21][19] = 4'hA;
    SS13[22][19] = 4'hA;
    SS13[23][19] = 4'hA;
    SS13[24][19] = 4'hA;
    SS13[25][19] = 4'hD;
    SS13[26][19] = 4'hD;
    SS13[27][19] = 4'hC;
    SS13[28][19] = 4'hC;
    SS13[29][19] = 4'hD;
    SS13[30][19] = 4'hD;
    SS13[31][19] = 4'hD;
    SS13[32][19] = 4'hD;
    SS13[33][19] = 4'hD;
    SS13[34][19] = 4'hD;
    SS13[35][19] = 4'hD;
    SS13[36][19] = 4'hD;
    SS13[37][19] = 4'hD;
    SS13[38][19] = 4'h3;
    SS13[39][19] = 4'h3;
    SS13[40][19] = 4'h3;
    SS13[41][19] = 4'h0;
    SS13[42][19] = 4'h0;
    SS13[43][19] = 4'hD;
    SS13[44][19] = 4'hD;
    SS13[45][19] = 4'h0;
    SS13[46][19] = 4'h0;
    SS13[47][19] = 4'h0;
    SS13[0][20] = 4'h0;
    SS13[1][20] = 4'h0;
    SS13[2][20] = 4'h0;
    SS13[3][20] = 4'h0;
    SS13[4][20] = 4'h0;
    SS13[5][20] = 4'h0;
    SS13[6][20] = 4'h0;
    SS13[7][20] = 4'h0;
    SS13[8][20] = 4'h0;
    SS13[9][20] = 4'h0;
    SS13[10][20] = 4'h0;
    SS13[11][20] = 4'h0;
    SS13[12][20] = 4'h0;
    SS13[13][20] = 4'h0;
    SS13[14][20] = 4'h0;
    SS13[15][20] = 4'h0;
    SS13[16][20] = 4'hC;
    SS13[17][20] = 4'hD;
    SS13[18][20] = 4'hD;
    SS13[19][20] = 4'hA;
    SS13[20][20] = 4'hA;
    SS13[21][20] = 4'hA;
    SS13[22][20] = 4'hA;
    SS13[23][20] = 4'hA;
    SS13[24][20] = 4'hA;
    SS13[25][20] = 4'hD;
    SS13[26][20] = 4'hC;
    SS13[27][20] = 4'hC;
    SS13[28][20] = 4'hC;
    SS13[29][20] = 4'hD;
    SS13[30][20] = 4'hD;
    SS13[31][20] = 4'hD;
    SS13[32][20] = 4'hD;
    SS13[33][20] = 4'hD;
    SS13[34][20] = 4'hD;
    SS13[35][20] = 4'hD;
    SS13[36][20] = 4'hD;
    SS13[37][20] = 4'hD;
    SS13[38][20] = 4'hD;
    SS13[39][20] = 4'h3;
    SS13[40][20] = 4'hD;
    SS13[41][20] = 4'hD;
    SS13[42][20] = 4'hD;
    SS13[43][20] = 4'hD;
    SS13[44][20] = 4'hD;
    SS13[45][20] = 4'h0;
    SS13[46][20] = 4'h0;
    SS13[47][20] = 4'h0;
    SS13[0][21] = 4'h0;
    SS13[1][21] = 4'h0;
    SS13[2][21] = 4'h0;
    SS13[3][21] = 4'h0;
    SS13[4][21] = 4'h0;
    SS13[5][21] = 4'h0;
    SS13[6][21] = 4'h0;
    SS13[7][21] = 4'h0;
    SS13[8][21] = 4'h0;
    SS13[9][21] = 4'h0;
    SS13[10][21] = 4'h0;
    SS13[11][21] = 4'h0;
    SS13[12][21] = 4'h0;
    SS13[13][21] = 4'h0;
    SS13[14][21] = 4'hF;
    SS13[15][21] = 4'hD;
    SS13[16][21] = 4'hD;
    SS13[17][21] = 4'hD;
    SS13[18][21] = 4'hD;
    SS13[19][21] = 4'hD;
    SS13[20][21] = 4'hA;
    SS13[21][21] = 4'hA;
    SS13[22][21] = 4'hD;
    SS13[23][21] = 4'hD;
    SS13[24][21] = 4'hD;
    SS13[25][21] = 4'hD;
    SS13[26][21] = 4'hC;
    SS13[27][21] = 4'hC;
    SS13[28][21] = 4'hC;
    SS13[29][21] = 4'hD;
    SS13[30][21] = 4'hE;
    SS13[31][21] = 4'hE;
    SS13[32][21] = 4'hE;
    SS13[33][21] = 4'hD;
    SS13[34][21] = 4'hD;
    SS13[35][21] = 4'hD;
    SS13[36][21] = 4'hD;
    SS13[37][21] = 4'hD;
    SS13[38][21] = 4'hE;
    SS13[39][21] = 4'hD;
    SS13[40][21] = 4'hD;
    SS13[41][21] = 4'hD;
    SS13[42][21] = 4'hD;
    SS13[43][21] = 4'hD;
    SS13[44][21] = 4'hD;
    SS13[45][21] = 4'hE;
    SS13[46][21] = 4'hD;
    SS13[47][21] = 4'hD;
    SS13[0][22] = 4'h0;
    SS13[1][22] = 4'h0;
    SS13[2][22] = 4'h0;
    SS13[3][22] = 4'h0;
    SS13[4][22] = 4'h0;
    SS13[5][22] = 4'h0;
    SS13[6][22] = 4'h0;
    SS13[7][22] = 4'h0;
    SS13[8][22] = 4'h0;
    SS13[9][22] = 4'h0;
    SS13[10][22] = 4'h0;
    SS13[11][22] = 4'h0;
    SS13[12][22] = 4'h3;
    SS13[13][22] = 4'h3;
    SS13[14][22] = 4'hD;
    SS13[15][22] = 4'hD;
    SS13[16][22] = 4'hD;
    SS13[17][22] = 4'hD;
    SS13[18][22] = 4'hD;
    SS13[19][22] = 4'hD;
    SS13[20][22] = 4'hD;
    SS13[21][22] = 4'hD;
    SS13[22][22] = 4'hD;
    SS13[23][22] = 4'hD;
    SS13[24][22] = 4'hD;
    SS13[25][22] = 4'hD;
    SS13[26][22] = 4'hD;
    SS13[27][22] = 4'hC;
    SS13[28][22] = 4'hC;
    SS13[29][22] = 4'hC;
    SS13[30][22] = 4'hE;
    SS13[31][22] = 4'hE;
    SS13[32][22] = 4'hE;
    SS13[33][22] = 4'hD;
    SS13[34][22] = 4'hD;
    SS13[35][22] = 4'hE;
    SS13[36][22] = 4'hE;
    SS13[37][22] = 4'hE;
    SS13[38][22] = 4'hE;
    SS13[39][22] = 4'hD;
    SS13[40][22] = 4'hD;
    SS13[41][22] = 4'hD;
    SS13[42][22] = 4'hD;
    SS13[43][22] = 4'hD;
    SS13[44][22] = 4'hD;
    SS13[45][22] = 4'hD;
    SS13[46][22] = 4'hD;
    SS13[47][22] = 4'hD;
    SS13[0][23] = 4'h0;
    SS13[1][23] = 4'h0;
    SS13[2][23] = 4'h0;
    SS13[3][23] = 4'h0;
    SS13[4][23] = 4'h0;
    SS13[5][23] = 4'h0;
    SS13[6][23] = 4'h0;
    SS13[7][23] = 4'h0;
    SS13[8][23] = 4'h0;
    SS13[9][23] = 4'h0;
    SS13[10][23] = 4'h0;
    SS13[11][23] = 4'h3;
    SS13[12][23] = 4'h3;
    SS13[13][23] = 4'h3;
    SS13[14][23] = 4'hD;
    SS13[15][23] = 4'hD;
    SS13[16][23] = 4'hD;
    SS13[17][23] = 4'hC;
    SS13[18][23] = 4'hC;
    SS13[19][23] = 4'hC;
    SS13[20][23] = 4'hC;
    SS13[21][23] = 4'hD;
    SS13[22][23] = 4'hD;
    SS13[23][23] = 4'hD;
    SS13[24][23] = 4'hD;
    SS13[25][23] = 4'hC;
    SS13[26][23] = 4'hC;
    SS13[27][23] = 4'hC;
    SS13[28][23] = 4'hC;
    SS13[29][23] = 4'hC;
    SS13[30][23] = 4'hE;
    SS13[31][23] = 4'hE;
    SS13[32][23] = 4'hE;
    SS13[33][23] = 4'hE;
    SS13[34][23] = 4'hE;
    SS13[35][23] = 4'hE;
    SS13[36][23] = 4'hE;
    SS13[37][23] = 4'hE;
    SS13[38][23] = 4'hE;
    SS13[39][23] = 4'hE;
    SS13[40][23] = 4'hD;
    SS13[41][23] = 4'hE;
    SS13[42][23] = 4'hE;
    SS13[43][23] = 4'hD;
    SS13[44][23] = 4'hD;
    SS13[45][23] = 4'hD;
    SS13[46][23] = 4'hD;
    SS13[47][23] = 4'hD;
    SS13[0][24] = 4'h0;
    SS13[1][24] = 4'h0;
    SS13[2][24] = 4'h0;
    SS13[3][24] = 4'h0;
    SS13[4][24] = 4'h0;
    SS13[5][24] = 4'h0;
    SS13[6][24] = 4'h0;
    SS13[7][24] = 4'h0;
    SS13[8][24] = 4'h0;
    SS13[9][24] = 4'h0;
    SS13[10][24] = 4'h0;
    SS13[11][24] = 4'h3;
    SS13[12][24] = 4'h3;
    SS13[13][24] = 4'h3;
    SS13[14][24] = 4'h3;
    SS13[15][24] = 4'hD;
    SS13[16][24] = 4'hD;
    SS13[17][24] = 4'hD;
    SS13[18][24] = 4'hC;
    SS13[19][24] = 4'hC;
    SS13[20][24] = 4'hC;
    SS13[21][24] = 4'hD;
    SS13[22][24] = 4'hD;
    SS13[23][24] = 4'hC;
    SS13[24][24] = 4'hC;
    SS13[25][24] = 4'hC;
    SS13[26][24] = 4'hC;
    SS13[27][24] = 4'hC;
    SS13[28][24] = 4'hC;
    SS13[29][24] = 4'hC;
    SS13[30][24] = 4'hC;
    SS13[31][24] = 4'hC;
    SS13[32][24] = 4'hC;
    SS13[33][24] = 4'hC;
    SS13[34][24] = 4'hE;
    SS13[35][24] = 4'hE;
    SS13[36][24] = 4'hE;
    SS13[37][24] = 4'hE;
    SS13[38][24] = 4'hE;
    SS13[39][24] = 4'hE;
    SS13[40][24] = 4'hE;
    SS13[41][24] = 4'hE;
    SS13[42][24] = 4'hE;
    SS13[43][24] = 4'hD;
    SS13[44][24] = 4'hD;
    SS13[45][24] = 4'hD;
    SS13[46][24] = 4'h0;
    SS13[47][24] = 4'h0;
    SS13[0][25] = 4'h0;
    SS13[1][25] = 4'h0;
    SS13[2][25] = 4'h0;
    SS13[3][25] = 4'h0;
    SS13[4][25] = 4'h0;
    SS13[5][25] = 4'h0;
    SS13[6][25] = 4'h0;
    SS13[7][25] = 4'h0;
    SS13[8][25] = 4'h0;
    SS13[9][25] = 4'h0;
    SS13[10][25] = 4'h0;
    SS13[11][25] = 4'h0;
    SS13[12][25] = 4'h3;
    SS13[13][25] = 4'hD;
    SS13[14][25] = 4'hD;
    SS13[15][25] = 4'hD;
    SS13[16][25] = 4'hD;
    SS13[17][25] = 4'hD;
    SS13[18][25] = 4'hC;
    SS13[19][25] = 4'hC;
    SS13[20][25] = 4'hC;
    SS13[21][25] = 4'hC;
    SS13[22][25] = 4'hC;
    SS13[23][25] = 4'hC;
    SS13[24][25] = 4'hC;
    SS13[25][25] = 4'hC;
    SS13[26][25] = 4'hC;
    SS13[27][25] = 4'hC;
    SS13[28][25] = 4'hC;
    SS13[29][25] = 4'hC;
    SS13[30][25] = 4'hC;
    SS13[31][25] = 4'hC;
    SS13[32][25] = 4'hC;
    SS13[33][25] = 4'hC;
    SS13[34][25] = 4'hE;
    SS13[35][25] = 4'hE;
    SS13[36][25] = 4'hC;
    SS13[37][25] = 4'hE;
    SS13[38][25] = 4'hE;
    SS13[39][25] = 4'hE;
    SS13[40][25] = 4'hE;
    SS13[41][25] = 4'hE;
    SS13[42][25] = 4'hE;
    SS13[43][25] = 4'hE;
    SS13[44][25] = 4'h0;
    SS13[45][25] = 4'h0;
    SS13[46][25] = 4'h0;
    SS13[47][25] = 4'h0;
    SS13[0][26] = 4'h0;
    SS13[1][26] = 4'h0;
    SS13[2][26] = 4'h0;
    SS13[3][26] = 4'h0;
    SS13[4][26] = 4'h0;
    SS13[5][26] = 4'h0;
    SS13[6][26] = 4'h0;
    SS13[7][26] = 4'h0;
    SS13[8][26] = 4'h0;
    SS13[9][26] = 4'h0;
    SS13[10][26] = 4'h0;
    SS13[11][26] = 4'h0;
    SS13[12][26] = 4'hD;
    SS13[13][26] = 4'hD;
    SS13[14][26] = 4'hD;
    SS13[15][26] = 4'hD;
    SS13[16][26] = 4'hD;
    SS13[17][26] = 4'hD;
    SS13[18][26] = 4'hE;
    SS13[19][26] = 4'hC;
    SS13[20][26] = 4'hC;
    SS13[21][26] = 4'hC;
    SS13[22][26] = 4'hC;
    SS13[23][26] = 4'hC;
    SS13[24][26] = 4'hC;
    SS13[25][26] = 4'hC;
    SS13[26][26] = 4'hD;
    SS13[27][26] = 4'hD;
    SS13[28][26] = 4'hC;
    SS13[29][26] = 4'hC;
    SS13[30][26] = 4'hC;
    SS13[31][26] = 4'hC;
    SS13[32][26] = 4'hC;
    SS13[33][26] = 4'hC;
    SS13[34][26] = 4'hC;
    SS13[35][26] = 4'hC;
    SS13[36][26] = 4'hC;
    SS13[37][26] = 4'hC;
    SS13[38][26] = 4'hE;
    SS13[39][26] = 4'hE;
    SS13[40][26] = 4'hE;
    SS13[41][26] = 4'h0;
    SS13[42][26] = 4'h0;
    SS13[43][26] = 4'h0;
    SS13[44][26] = 4'h0;
    SS13[45][26] = 4'h0;
    SS13[46][26] = 4'h0;
    SS13[47][26] = 4'h0;
    SS13[0][27] = 4'h0;
    SS13[1][27] = 4'h0;
    SS13[2][27] = 4'h0;
    SS13[3][27] = 4'h0;
    SS13[4][27] = 4'h0;
    SS13[5][27] = 4'h0;
    SS13[6][27] = 4'h0;
    SS13[7][27] = 4'h0;
    SS13[8][27] = 4'h0;
    SS13[9][27] = 4'h0;
    SS13[10][27] = 4'h0;
    SS13[11][27] = 4'h0;
    SS13[12][27] = 4'h0;
    SS13[13][27] = 4'hD;
    SS13[14][27] = 4'hD;
    SS13[15][27] = 4'hD;
    SS13[16][27] = 4'hE;
    SS13[17][27] = 4'hE;
    SS13[18][27] = 4'hE;
    SS13[19][27] = 4'hC;
    SS13[20][27] = 4'hC;
    SS13[21][27] = 4'hC;
    SS13[22][27] = 4'hC;
    SS13[23][27] = 4'hD;
    SS13[24][27] = 4'hD;
    SS13[25][27] = 4'hD;
    SS13[26][27] = 4'hD;
    SS13[27][27] = 4'hD;
    SS13[28][27] = 4'hD;
    SS13[29][27] = 4'hC;
    SS13[30][27] = 4'hC;
    SS13[31][27] = 4'hC;
    SS13[32][27] = 4'hC;
    SS13[33][27] = 4'hC;
    SS13[34][27] = 4'hC;
    SS13[35][27] = 4'hC;
    SS13[36][27] = 4'hC;
    SS13[37][27] = 4'hC;
    SS13[38][27] = 4'hE;
    SS13[39][27] = 4'h0;
    SS13[40][27] = 4'h0;
    SS13[41][27] = 4'h0;
    SS13[42][27] = 4'h0;
    SS13[43][27] = 4'h0;
    SS13[44][27] = 4'h0;
    SS13[45][27] = 4'h0;
    SS13[46][27] = 4'h0;
    SS13[47][27] = 4'h0;
    SS13[0][28] = 4'h0;
    SS13[1][28] = 4'h0;
    SS13[2][28] = 4'h0;
    SS13[3][28] = 4'h0;
    SS13[4][28] = 4'h0;
    SS13[5][28] = 4'h0;
    SS13[6][28] = 4'h0;
    SS13[7][28] = 4'h0;
    SS13[8][28] = 4'h0;
    SS13[9][28] = 4'h0;
    SS13[10][28] = 4'h0;
    SS13[11][28] = 4'h0;
    SS13[12][28] = 4'h0;
    SS13[13][28] = 4'hD;
    SS13[14][28] = 4'hD;
    SS13[15][28] = 4'hD;
    SS13[16][28] = 4'hE;
    SS13[17][28] = 4'hE;
    SS13[18][28] = 4'hE;
    SS13[19][28] = 4'hC;
    SS13[20][28] = 4'hC;
    SS13[21][28] = 4'hC;
    SS13[22][28] = 4'hC;
    SS13[23][28] = 4'hD;
    SS13[24][28] = 4'hD;
    SS13[25][28] = 4'hD;
    SS13[26][28] = 4'hD;
    SS13[27][28] = 4'hD;
    SS13[28][28] = 4'hD;
    SS13[29][28] = 4'hC;
    SS13[30][28] = 4'hC;
    SS13[31][28] = 4'hC;
    SS13[32][28] = 4'hC;
    SS13[33][28] = 4'hC;
    SS13[34][28] = 4'hC;
    SS13[35][28] = 4'hC;
    SS13[36][28] = 4'hC;
    SS13[37][28] = 4'hC;
    SS13[38][28] = 4'hC;
    SS13[39][28] = 4'h0;
    SS13[40][28] = 4'h0;
    SS13[41][28] = 4'h0;
    SS13[42][28] = 4'h0;
    SS13[43][28] = 4'h0;
    SS13[44][28] = 4'h0;
    SS13[45][28] = 4'h0;
    SS13[46][28] = 4'h0;
    SS13[47][28] = 4'h0;
    SS13[0][29] = 4'h0;
    SS13[1][29] = 4'h0;
    SS13[2][29] = 4'h0;
    SS13[3][29] = 4'h0;
    SS13[4][29] = 4'h0;
    SS13[5][29] = 4'h0;
    SS13[6][29] = 4'h0;
    SS13[7][29] = 4'h0;
    SS13[8][29] = 4'h0;
    SS13[9][29] = 4'h0;
    SS13[10][29] = 4'h0;
    SS13[11][29] = 4'hD;
    SS13[12][29] = 4'hD;
    SS13[13][29] = 4'hD;
    SS13[14][29] = 4'hD;
    SS13[15][29] = 4'hD;
    SS13[16][29] = 4'hD;
    SS13[17][29] = 4'hE;
    SS13[18][29] = 4'hC;
    SS13[19][29] = 4'hC;
    SS13[20][29] = 4'hC;
    SS13[21][29] = 4'hC;
    SS13[22][29] = 4'hC;
    SS13[23][29] = 4'hD;
    SS13[24][29] = 4'hD;
    SS13[25][29] = 4'hD;
    SS13[26][29] = 4'hE;
    SS13[27][29] = 4'hE;
    SS13[28][29] = 4'hE;
    SS13[29][29] = 4'hC;
    SS13[30][29] = 4'hC;
    SS13[31][29] = 4'hC;
    SS13[32][29] = 4'hC;
    SS13[33][29] = 4'hC;
    SS13[34][29] = 4'hC;
    SS13[35][29] = 4'hC;
    SS13[36][29] = 4'hC;
    SS13[37][29] = 4'hC;
    SS13[38][29] = 4'hC;
    SS13[39][29] = 4'h0;
    SS13[40][29] = 4'h0;
    SS13[41][29] = 4'h0;
    SS13[42][29] = 4'h0;
    SS13[43][29] = 4'h0;
    SS13[44][29] = 4'h0;
    SS13[45][29] = 4'h0;
    SS13[46][29] = 4'h0;
    SS13[47][29] = 4'h0;
    SS13[0][30] = 4'h0;
    SS13[1][30] = 4'h0;
    SS13[2][30] = 4'h0;
    SS13[3][30] = 4'h0;
    SS13[4][30] = 4'h0;
    SS13[5][30] = 4'h0;
    SS13[6][30] = 4'h0;
    SS13[7][30] = 4'h0;
    SS13[8][30] = 4'h3;
    SS13[9][30] = 4'h3;
    SS13[10][30] = 4'h3;
    SS13[11][30] = 4'hD;
    SS13[12][30] = 4'hD;
    SS13[13][30] = 4'hD;
    SS13[14][30] = 4'hD;
    SS13[15][30] = 4'hD;
    SS13[16][30] = 4'hE;
    SS13[17][30] = 4'hC;
    SS13[18][30] = 4'hC;
    SS13[19][30] = 4'hC;
    SS13[20][30] = 4'hC;
    SS13[21][30] = 4'hC;
    SS13[22][30] = 4'hC;
    SS13[23][30] = 4'hD;
    SS13[24][30] = 4'hE;
    SS13[25][30] = 4'hE;
    SS13[26][30] = 4'hE;
    SS13[27][30] = 4'hE;
    SS13[28][30] = 4'hE;
    SS13[29][30] = 4'hE;
    SS13[30][30] = 4'hC;
    SS13[31][30] = 4'hC;
    SS13[32][30] = 4'hD;
    SS13[33][30] = 4'hC;
    SS13[34][30] = 4'hC;
    SS13[35][30] = 4'hC;
    SS13[36][30] = 4'hC;
    SS13[37][30] = 4'hC;
    SS13[38][30] = 4'hC;
    SS13[39][30] = 4'hC;
    SS13[40][30] = 4'h0;
    SS13[41][30] = 4'h0;
    SS13[42][30] = 4'h0;
    SS13[43][30] = 4'h0;
    SS13[44][30] = 4'h0;
    SS13[45][30] = 4'h0;
    SS13[46][30] = 4'h0;
    SS13[47][30] = 4'h0;
    SS13[0][31] = 4'h0;
    SS13[1][31] = 4'h0;
    SS13[2][31] = 4'h0;
    SS13[3][31] = 4'h0;
    SS13[4][31] = 4'h0;
    SS13[5][31] = 4'h0;
    SS13[6][31] = 4'h0;
    SS13[7][31] = 4'h0;
    SS13[8][31] = 4'h3;
    SS13[9][31] = 4'h3;
    SS13[10][31] = 4'h3;
    SS13[11][31] = 4'hD;
    SS13[12][31] = 4'hD;
    SS13[13][31] = 4'hD;
    SS13[14][31] = 4'hE;
    SS13[15][31] = 4'hE;
    SS13[16][31] = 4'hE;
    SS13[17][31] = 4'hC;
    SS13[18][31] = 4'hC;
    SS13[19][31] = 4'hC;
    SS13[20][31] = 4'hC;
    SS13[21][31] = 4'hC;
    SS13[22][31] = 4'hC;
    SS13[23][31] = 4'hC;
    SS13[24][31] = 4'hE;
    SS13[25][31] = 4'hE;
    SS13[26][31] = 4'hE;
    SS13[27][31] = 4'hE;
    SS13[28][31] = 4'hE;
    SS13[29][31] = 4'hE;
    SS13[30][31] = 4'hD;
    SS13[31][31] = 4'hD;
    SS13[32][31] = 4'hD;
    SS13[33][31] = 4'hD;
    SS13[34][31] = 4'hC;
    SS13[35][31] = 4'hC;
    SS13[36][31] = 4'hC;
    SS13[37][31] = 4'hC;
    SS13[38][31] = 4'hC;
    SS13[39][31] = 4'hC;
    SS13[40][31] = 4'h0;
    SS13[41][31] = 4'h0;
    SS13[42][31] = 4'h0;
    SS13[43][31] = 4'h0;
    SS13[44][31] = 4'h0;
    SS13[45][31] = 4'h0;
    SS13[46][31] = 4'h0;
    SS13[47][31] = 4'h0;
    SS13[0][32] = 4'h0;
    SS13[1][32] = 4'h0;
    SS13[2][32] = 4'h0;
    SS13[3][32] = 4'h0;
    SS13[4][32] = 4'h0;
    SS13[5][32] = 4'h0;
    SS13[6][32] = 4'h0;
    SS13[7][32] = 4'h0;
    SS13[8][32] = 4'h3;
    SS13[9][32] = 4'h3;
    SS13[10][32] = 4'h3;
    SS13[11][32] = 4'hE;
    SS13[12][32] = 4'hE;
    SS13[13][32] = 4'hE;
    SS13[14][32] = 4'hE;
    SS13[15][32] = 4'hE;
    SS13[16][32] = 4'hE;
    SS13[17][32] = 4'hE;
    SS13[18][32] = 4'hC;
    SS13[19][32] = 4'hC;
    SS13[20][32] = 4'hC;
    SS13[21][32] = 4'hC;
    SS13[22][32] = 4'hC;
    SS13[23][32] = 4'hC;
    SS13[24][32] = 4'hE;
    SS13[25][32] = 4'hE;
    SS13[26][32] = 4'hE;
    SS13[27][32] = 4'hE;
    SS13[28][32] = 4'hE;
    SS13[29][32] = 4'hE;
    SS13[30][32] = 4'hE;
    SS13[31][32] = 4'hD;
    SS13[32][32] = 4'hD;
    SS13[33][32] = 4'hD;
    SS13[34][32] = 4'hD;
    SS13[35][32] = 4'hD;
    SS13[36][32] = 4'hD;
    SS13[37][32] = 4'hC;
    SS13[38][32] = 4'hC;
    SS13[39][32] = 4'hC;
    SS13[40][32] = 4'h0;
    SS13[41][32] = 4'h0;
    SS13[42][32] = 4'hC;
    SS13[43][32] = 4'hC;
    SS13[44][32] = 4'h0;
    SS13[45][32] = 4'h0;
    SS13[46][32] = 4'h0;
    SS13[47][32] = 4'h0;
    SS13[0][33] = 4'h0;
    SS13[1][33] = 4'h0;
    SS13[2][33] = 4'h0;
    SS13[3][33] = 4'h0;
    SS13[4][33] = 4'h0;
    SS13[5][33] = 4'h0;
    SS13[6][33] = 4'h0;
    SS13[7][33] = 4'h0;
    SS13[8][33] = 4'h0;
    SS13[9][33] = 4'hD;
    SS13[10][33] = 4'hD;
    SS13[11][33] = 4'hD;
    SS13[12][33] = 4'hE;
    SS13[13][33] = 4'hE;
    SS13[14][33] = 4'hE;
    SS13[15][33] = 4'hE;
    SS13[16][33] = 4'hE;
    SS13[17][33] = 4'hC;
    SS13[18][33] = 4'hC;
    SS13[19][33] = 4'hC;
    SS13[20][33] = 4'hC;
    SS13[21][33] = 4'hC;
    SS13[22][33] = 4'hC;
    SS13[23][33] = 4'hC;
    SS13[24][33] = 4'hD;
    SS13[25][33] = 4'hE;
    SS13[26][33] = 4'hE;
    SS13[27][33] = 4'hE;
    SS13[28][33] = 4'hE;
    SS13[29][33] = 4'hE;
    SS13[30][33] = 4'hE;
    SS13[31][33] = 4'hD;
    SS13[32][33] = 4'hE;
    SS13[33][33] = 4'hE;
    SS13[34][33] = 4'hD;
    SS13[35][33] = 4'hD;
    SS13[36][33] = 4'hD;
    SS13[37][33] = 4'hD;
    SS13[38][33] = 4'hC;
    SS13[39][33] = 4'hC;
    SS13[40][33] = 4'hC;
    SS13[41][33] = 4'hC;
    SS13[42][33] = 4'hC;
    SS13[43][33] = 4'hC;
    SS13[44][33] = 4'h0;
    SS13[45][33] = 4'h0;
    SS13[46][33] = 4'h0;
    SS13[47][33] = 4'h0;
    SS13[0][34] = 4'h0;
    SS13[1][34] = 4'h0;
    SS13[2][34] = 4'h0;
    SS13[3][34] = 4'h0;
    SS13[4][34] = 4'h0;
    SS13[5][34] = 4'h0;
    SS13[6][34] = 4'hD;
    SS13[7][34] = 4'hD;
    SS13[8][34] = 4'hD;
    SS13[9][34] = 4'hD;
    SS13[10][34] = 4'hD;
    SS13[11][34] = 4'hD;
    SS13[12][34] = 4'hE;
    SS13[13][34] = 4'hE;
    SS13[14][34] = 4'hE;
    SS13[15][34] = 4'hE;
    SS13[16][34] = 4'hC;
    SS13[17][34] = 4'hC;
    SS13[18][34] = 4'hC;
    SS13[19][34] = 4'hC;
    SS13[20][34] = 4'hC;
    SS13[21][34] = 4'hC;
    SS13[22][34] = 4'hD;
    SS13[23][34] = 4'hD;
    SS13[24][34] = 4'hD;
    SS13[25][34] = 4'hE;
    SS13[26][34] = 4'hE;
    SS13[27][34] = 4'hE;
    SS13[28][34] = 4'hE;
    SS13[29][34] = 4'hE;
    SS13[30][34] = 4'h0;
    SS13[31][34] = 4'h0;
    SS13[32][34] = 4'hE;
    SS13[33][34] = 4'hE;
    SS13[34][34] = 4'hE;
    SS13[35][34] = 4'hD;
    SS13[36][34] = 4'hD;
    SS13[37][34] = 4'hE;
    SS13[38][34] = 4'hC;
    SS13[39][34] = 4'hC;
    SS13[40][34] = 4'hC;
    SS13[41][34] = 4'hC;
    SS13[42][34] = 4'hC;
    SS13[43][34] = 4'hC;
    SS13[44][34] = 4'h0;
    SS13[45][34] = 4'h0;
    SS13[46][34] = 4'h0;
    SS13[47][34] = 4'h0;
    SS13[0][35] = 4'h0;
    SS13[1][35] = 4'h0;
    SS13[2][35] = 4'h0;
    SS13[3][35] = 4'h0;
    SS13[4][35] = 4'h0;
    SS13[5][35] = 4'h0;
    SS13[6][35] = 4'hD;
    SS13[7][35] = 4'hD;
    SS13[8][35] = 4'hD;
    SS13[9][35] = 4'hD;
    SS13[10][35] = 4'hD;
    SS13[11][35] = 4'hD;
    SS13[12][35] = 4'hE;
    SS13[13][35] = 4'hE;
    SS13[14][35] = 4'hE;
    SS13[15][35] = 4'hE;
    SS13[16][35] = 4'hC;
    SS13[17][35] = 4'hC;
    SS13[18][35] = 4'hC;
    SS13[19][35] = 4'hC;
    SS13[20][35] = 4'hC;
    SS13[21][35] = 4'hC;
    SS13[22][35] = 4'hD;
    SS13[23][35] = 4'hD;
    SS13[24][35] = 4'hD;
    SS13[25][35] = 4'hD;
    SS13[26][35] = 4'hE;
    SS13[27][35] = 4'h0;
    SS13[28][35] = 4'h0;
    SS13[29][35] = 4'h0;
    SS13[30][35] = 4'h0;
    SS13[31][35] = 4'h0;
    SS13[32][35] = 4'hE;
    SS13[33][35] = 4'hE;
    SS13[34][35] = 4'hE;
    SS13[35][35] = 4'hE;
    SS13[36][35] = 4'hE;
    SS13[37][35] = 4'hE;
    SS13[38][35] = 4'hC;
    SS13[39][35] = 4'hC;
    SS13[40][35] = 4'hC;
    SS13[41][35] = 4'hC;
    SS13[42][35] = 4'hC;
    SS13[43][35] = 4'hC;
    SS13[44][35] = 4'hC;
    SS13[45][35] = 4'h0;
    SS13[46][35] = 4'h0;
    SS13[47][35] = 4'h0;
    SS13[0][36] = 4'h0;
    SS13[1][36] = 4'h0;
    SS13[2][36] = 4'h0;
    SS13[3][36] = 4'h0;
    SS13[4][36] = 4'h0;
    SS13[5][36] = 4'h0;
    SS13[6][36] = 4'h0;
    SS13[7][36] = 4'hD;
    SS13[8][36] = 4'hD;
    SS13[9][36] = 4'hD;
    SS13[10][36] = 4'hE;
    SS13[11][36] = 4'hE;
    SS13[12][36] = 4'hE;
    SS13[13][36] = 4'hE;
    SS13[14][36] = 4'hE;
    SS13[15][36] = 4'hE;
    SS13[16][36] = 4'hC;
    SS13[17][36] = 4'hC;
    SS13[18][36] = 4'hC;
    SS13[19][36] = 4'hC;
    SS13[20][36] = 4'hC;
    SS13[21][36] = 4'hC;
    SS13[22][36] = 4'hC;
    SS13[23][36] = 4'hD;
    SS13[24][36] = 4'hD;
    SS13[25][36] = 4'hE;
    SS13[26][36] = 4'h0;
    SS13[27][36] = 4'h0;
    SS13[28][36] = 4'h0;
    SS13[29][36] = 4'h0;
    SS13[30][36] = 4'h0;
    SS13[31][36] = 4'h0;
    SS13[32][36] = 4'hE;
    SS13[33][36] = 4'h0;
    SS13[34][36] = 4'h0;
    SS13[35][36] = 4'h0;
    SS13[36][36] = 4'hE;
    SS13[37][36] = 4'hE;
    SS13[38][36] = 4'hE;
    SS13[39][36] = 4'hC;
    SS13[40][36] = 4'hD;
    SS13[41][36] = 4'hD;
    SS13[42][36] = 4'hC;
    SS13[43][36] = 4'hC;
    SS13[44][36] = 4'hC;
    SS13[45][36] = 4'h0;
    SS13[46][36] = 4'h0;
    SS13[47][36] = 4'h0;
    SS13[0][37] = 4'h0;
    SS13[1][37] = 4'h0;
    SS13[2][37] = 4'h0;
    SS13[3][37] = 4'h0;
    SS13[4][37] = 4'h0;
    SS13[5][37] = 4'h0;
    SS13[6][37] = 4'h0;
    SS13[7][37] = 4'hD;
    SS13[8][37] = 4'hD;
    SS13[9][37] = 4'hD;
    SS13[10][37] = 4'hE;
    SS13[11][37] = 4'hE;
    SS13[12][37] = 4'hE;
    SS13[13][37] = 4'hE;
    SS13[14][37] = 4'hE;
    SS13[15][37] = 4'h0;
    SS13[16][37] = 4'h0;
    SS13[17][37] = 4'hC;
    SS13[18][37] = 4'hC;
    SS13[19][37] = 4'hC;
    SS13[20][37] = 4'hC;
    SS13[21][37] = 4'hC;
    SS13[22][37] = 4'hD;
    SS13[23][37] = 4'hE;
    SS13[24][37] = 4'hE;
    SS13[25][37] = 4'hE;
    SS13[26][37] = 4'h0;
    SS13[27][37] = 4'h0;
    SS13[28][37] = 4'h0;
    SS13[29][37] = 4'h0;
    SS13[30][37] = 4'h0;
    SS13[31][37] = 4'h0;
    SS13[32][37] = 4'h0;
    SS13[33][37] = 4'h0;
    SS13[34][37] = 4'h0;
    SS13[35][37] = 4'h0;
    SS13[36][37] = 4'hE;
    SS13[37][37] = 4'hE;
    SS13[38][37] = 4'h0;
    SS13[39][37] = 4'hD;
    SS13[40][37] = 4'hD;
    SS13[41][37] = 4'hD;
    SS13[42][37] = 4'hC;
    SS13[43][37] = 4'hC;
    SS13[44][37] = 4'hC;
    SS13[45][37] = 4'hC;
    SS13[46][37] = 4'h0;
    SS13[47][37] = 4'h0;
    SS13[0][38] = 4'h0;
    SS13[1][38] = 4'h0;
    SS13[2][38] = 4'h0;
    SS13[3][38] = 4'h0;
    SS13[4][38] = 4'hD;
    SS13[5][38] = 4'hD;
    SS13[6][38] = 4'hD;
    SS13[7][38] = 4'hD;
    SS13[8][38] = 4'hD;
    SS13[9][38] = 4'hD;
    SS13[10][38] = 4'hD;
    SS13[11][38] = 4'hE;
    SS13[12][38] = 4'h0;
    SS13[13][38] = 4'h0;
    SS13[14][38] = 4'h0;
    SS13[15][38] = 4'h0;
    SS13[16][38] = 4'h0;
    SS13[17][38] = 4'hC;
    SS13[18][38] = 4'hC;
    SS13[19][38] = 4'hC;
    SS13[20][38] = 4'hD;
    SS13[21][38] = 4'hD;
    SS13[22][38] = 4'hD;
    SS13[23][38] = 4'hD;
    SS13[24][38] = 4'hE;
    SS13[25][38] = 4'hE;
    SS13[26][38] = 4'hE;
    SS13[27][38] = 4'h0;
    SS13[28][38] = 4'h0;
    SS13[29][38] = 4'h0;
    SS13[30][38] = 4'h0;
    SS13[31][38] = 4'h0;
    SS13[32][38] = 4'h0;
    SS13[33][38] = 4'h0;
    SS13[34][38] = 4'h0;
    SS13[35][38] = 4'h0;
    SS13[36][38] = 4'h0;
    SS13[37][38] = 4'h0;
    SS13[38][38] = 4'h0;
    SS13[39][38] = 4'h0;
    SS13[40][38] = 4'hD;
    SS13[41][38] = 4'hD;
    SS13[42][38] = 4'hD;
    SS13[43][38] = 4'hD;
    SS13[44][38] = 4'hD;
    SS13[45][38] = 4'hD;
    SS13[46][38] = 4'h0;
    SS13[47][38] = 4'h0;
    SS13[0][39] = 4'h0;
    SS13[1][39] = 4'h0;
    SS13[2][39] = 4'h0;
    SS13[3][39] = 4'h0;
    SS13[4][39] = 4'h0;
    SS13[5][39] = 4'hD;
    SS13[6][39] = 4'hD;
    SS13[7][39] = 4'hD;
    SS13[8][39] = 4'hD;
    SS13[9][39] = 4'hD;
    SS13[10][39] = 4'h0;
    SS13[11][39] = 4'h0;
    SS13[12][39] = 4'h0;
    SS13[13][39] = 4'h0;
    SS13[14][39] = 4'h0;
    SS13[15][39] = 4'h0;
    SS13[16][39] = 4'h0;
    SS13[17][39] = 4'h0;
    SS13[18][39] = 4'hC;
    SS13[19][39] = 4'hC;
    SS13[20][39] = 4'hC;
    SS13[21][39] = 4'hD;
    SS13[22][39] = 4'hD;
    SS13[23][39] = 4'hD;
    SS13[24][39] = 4'hE;
    SS13[25][39] = 4'h0;
    SS13[26][39] = 4'h0;
    SS13[27][39] = 4'h0;
    SS13[28][39] = 4'h0;
    SS13[29][39] = 4'h0;
    SS13[30][39] = 4'h0;
    SS13[31][39] = 4'h0;
    SS13[32][39] = 4'h0;
    SS13[33][39] = 4'h0;
    SS13[34][39] = 4'h0;
    SS13[35][39] = 4'h0;
    SS13[36][39] = 4'h0;
    SS13[37][39] = 4'h0;
    SS13[38][39] = 4'h0;
    SS13[39][39] = 4'h0;
    SS13[40][39] = 4'hD;
    SS13[41][39] = 4'h0;
    SS13[42][39] = 4'h0;
    SS13[43][39] = 4'hD;
    SS13[44][39] = 4'hD;
    SS13[45][39] = 4'hD;
    SS13[46][39] = 4'h0;
    SS13[47][39] = 4'h0;
    SS13[0][40] = 4'h0;
    SS13[1][40] = 4'h0;
    SS13[2][40] = 4'h0;
    SS13[3][40] = 4'h0;
    SS13[4][40] = 4'h0;
    SS13[5][40] = 4'hD;
    SS13[6][40] = 4'hD;
    SS13[7][40] = 4'h0;
    SS13[8][40] = 4'h0;
    SS13[9][40] = 4'h0;
    SS13[10][40] = 4'h0;
    SS13[11][40] = 4'h0;
    SS13[12][40] = 4'h0;
    SS13[13][40] = 4'h0;
    SS13[14][40] = 4'h0;
    SS13[15][40] = 4'h0;
    SS13[16][40] = 4'h0;
    SS13[17][40] = 4'h0;
    SS13[18][40] = 4'hC;
    SS13[19][40] = 4'hC;
    SS13[20][40] = 4'hC;
    SS13[21][40] = 4'hD;
    SS13[22][40] = 4'hD;
    SS13[23][40] = 4'hE;
    SS13[24][40] = 4'h0;
    SS13[25][40] = 4'h0;
    SS13[26][40] = 4'h0;
    SS13[27][40] = 4'h0;
    SS13[28][40] = 4'h0;
    SS13[29][40] = 4'h0;
    SS13[30][40] = 4'h0;
    SS13[31][40] = 4'h0;
    SS13[32][40] = 4'h0;
    SS13[33][40] = 4'h0;
    SS13[34][40] = 4'h0;
    SS13[35][40] = 4'h0;
    SS13[36][40] = 4'h0;
    SS13[37][40] = 4'h0;
    SS13[38][40] = 4'h0;
    SS13[39][40] = 4'h0;
    SS13[40][40] = 4'h0;
    SS13[41][40] = 4'h0;
    SS13[42][40] = 4'h0;
    SS13[43][40] = 4'h0;
    SS13[44][40] = 4'hD;
    SS13[45][40] = 4'hD;
    SS13[46][40] = 4'h0;
    SS13[47][40] = 4'h0;
    SS13[0][41] = 4'h0;
    SS13[1][41] = 4'h0;
    SS13[2][41] = 4'h0;
    SS13[3][41] = 4'h0;
    SS13[4][41] = 4'h0;
    SS13[5][41] = 4'h0;
    SS13[6][41] = 4'h0;
    SS13[7][41] = 4'h0;
    SS13[8][41] = 4'h0;
    SS13[9][41] = 4'h0;
    SS13[10][41] = 4'h0;
    SS13[11][41] = 4'h0;
    SS13[12][41] = 4'h0;
    SS13[13][41] = 4'h0;
    SS13[14][41] = 4'h0;
    SS13[15][41] = 4'h0;
    SS13[16][41] = 4'h0;
    SS13[17][41] = 4'h0;
    SS13[18][41] = 4'hC;
    SS13[19][41] = 4'hC;
    SS13[20][41] = 4'hC;
    SS13[21][41] = 4'hC;
    SS13[22][41] = 4'hE;
    SS13[23][41] = 4'hE;
    SS13[24][41] = 4'hE;
    SS13[25][41] = 4'h0;
    SS13[26][41] = 4'h0;
    SS13[27][41] = 4'h0;
    SS13[28][41] = 4'h0;
    SS13[29][41] = 4'h0;
    SS13[30][41] = 4'h0;
    SS13[31][41] = 4'h0;
    SS13[32][41] = 4'h0;
    SS13[33][41] = 4'h0;
    SS13[34][41] = 4'h0;
    SS13[35][41] = 4'h0;
    SS13[36][41] = 4'h0;
    SS13[37][41] = 4'h0;
    SS13[38][41] = 4'h0;
    SS13[39][41] = 4'h0;
    SS13[40][41] = 4'h0;
    SS13[41][41] = 4'h0;
    SS13[42][41] = 4'h0;
    SS13[43][41] = 4'h0;
    SS13[44][41] = 4'h0;
    SS13[45][41] = 4'h0;
    SS13[46][41] = 4'h0;
    SS13[47][41] = 4'h0;
    SS13[0][42] = 4'h0;
    SS13[1][42] = 4'h0;
    SS13[2][42] = 4'h0;
    SS13[3][42] = 4'h0;
    SS13[4][42] = 4'h0;
    SS13[5][42] = 4'h0;
    SS13[6][42] = 4'h0;
    SS13[7][42] = 4'h0;
    SS13[8][42] = 4'h0;
    SS13[9][42] = 4'h0;
    SS13[10][42] = 4'h0;
    SS13[11][42] = 4'h0;
    SS13[12][42] = 4'h0;
    SS13[13][42] = 4'h0;
    SS13[14][42] = 4'h0;
    SS13[15][42] = 4'h0;
    SS13[16][42] = 4'h0;
    SS13[17][42] = 4'h0;
    SS13[18][42] = 4'hC;
    SS13[19][42] = 4'hC;
    SS13[20][42] = 4'hC;
    SS13[21][42] = 4'hC;
    SS13[22][42] = 4'hE;
    SS13[23][42] = 4'hE;
    SS13[24][42] = 4'hE;
    SS13[25][42] = 4'h0;
    SS13[26][42] = 4'h0;
    SS13[27][42] = 4'h0;
    SS13[28][42] = 4'h0;
    SS13[29][42] = 4'h0;
    SS13[30][42] = 4'h0;
    SS13[31][42] = 4'h0;
    SS13[32][42] = 4'h0;
    SS13[33][42] = 4'h0;
    SS13[34][42] = 4'h0;
    SS13[35][42] = 4'h0;
    SS13[36][42] = 4'h0;
    SS13[37][42] = 4'h0;
    SS13[38][42] = 4'h0;
    SS13[39][42] = 4'h0;
    SS13[40][42] = 4'h0;
    SS13[41][42] = 4'h0;
    SS13[42][42] = 4'h0;
    SS13[43][42] = 4'h0;
    SS13[44][42] = 4'h0;
    SS13[45][42] = 4'h0;
    SS13[46][42] = 4'h0;
    SS13[47][42] = 4'h0;
    SS13[0][43] = 4'h0;
    SS13[1][43] = 4'h0;
    SS13[2][43] = 4'h0;
    SS13[3][43] = 4'h0;
    SS13[4][43] = 4'h0;
    SS13[5][43] = 4'h0;
    SS13[6][43] = 4'h0;
    SS13[7][43] = 4'h0;
    SS13[8][43] = 4'h0;
    SS13[9][43] = 4'h0;
    SS13[10][43] = 4'h0;
    SS13[11][43] = 4'h0;
    SS13[12][43] = 4'h0;
    SS13[13][43] = 4'h0;
    SS13[14][43] = 4'h0;
    SS13[15][43] = 4'h0;
    SS13[16][43] = 4'hC;
    SS13[17][43] = 4'hC;
    SS13[18][43] = 4'hC;
    SS13[19][43] = 4'hC;
    SS13[20][43] = 4'hC;
    SS13[21][43] = 4'hC;
    SS13[22][43] = 4'hE;
    SS13[23][43] = 4'h0;
    SS13[24][43] = 4'h0;
    SS13[25][43] = 4'h0;
    SS13[26][43] = 4'h0;
    SS13[27][43] = 4'h0;
    SS13[28][43] = 4'h0;
    SS13[29][43] = 4'h0;
    SS13[30][43] = 4'h0;
    SS13[31][43] = 4'h0;
    SS13[32][43] = 4'h0;
    SS13[33][43] = 4'h0;
    SS13[34][43] = 4'h0;
    SS13[35][43] = 4'h0;
    SS13[36][43] = 4'h0;
    SS13[37][43] = 4'h0;
    SS13[38][43] = 4'h0;
    SS13[39][43] = 4'h0;
    SS13[40][43] = 4'h0;
    SS13[41][43] = 4'h0;
    SS13[42][43] = 4'h0;
    SS13[43][43] = 4'h0;
    SS13[44][43] = 4'h0;
    SS13[45][43] = 4'h0;
    SS13[46][43] = 4'h0;
    SS13[47][43] = 4'h0;
    SS13[0][44] = 4'h0;
    SS13[1][44] = 4'h0;
    SS13[2][44] = 4'h0;
    SS13[3][44] = 4'h0;
    SS13[4][44] = 4'h0;
    SS13[5][44] = 4'h0;
    SS13[6][44] = 4'h0;
    SS13[7][44] = 4'h0;
    SS13[8][44] = 4'h0;
    SS13[9][44] = 4'h0;
    SS13[10][44] = 4'h0;
    SS13[11][44] = 4'h0;
    SS13[12][44] = 4'h0;
    SS13[13][44] = 4'h0;
    SS13[14][44] = 4'h0;
    SS13[15][44] = 4'h0;
    SS13[16][44] = 4'hC;
    SS13[17][44] = 4'hC;
    SS13[18][44] = 4'hC;
    SS13[19][44] = 4'hC;
    SS13[20][44] = 4'hC;
    SS13[21][44] = 4'hD;
    SS13[22][44] = 4'hD;
    SS13[23][44] = 4'h0;
    SS13[24][44] = 4'h0;
    SS13[25][44] = 4'h0;
    SS13[26][44] = 4'h0;
    SS13[27][44] = 4'h0;
    SS13[28][44] = 4'h0;
    SS13[29][44] = 4'h0;
    SS13[30][44] = 4'h0;
    SS13[31][44] = 4'h0;
    SS13[32][44] = 4'h0;
    SS13[33][44] = 4'h0;
    SS13[34][44] = 4'h0;
    SS13[35][44] = 4'h0;
    SS13[36][44] = 4'h0;
    SS13[37][44] = 4'h0;
    SS13[38][44] = 4'h0;
    SS13[39][44] = 4'h0;
    SS13[40][44] = 4'h0;
    SS13[41][44] = 4'h0;
    SS13[42][44] = 4'h0;
    SS13[43][44] = 4'h0;
    SS13[44][44] = 4'h0;
    SS13[45][44] = 4'h0;
    SS13[46][44] = 4'h0;
    SS13[47][44] = 4'h0;
    SS13[0][45] = 4'h0;
    SS13[1][45] = 4'h0;
    SS13[2][45] = 4'h0;
    SS13[3][45] = 4'h0;
    SS13[4][45] = 4'h0;
    SS13[5][45] = 4'h0;
    SS13[6][45] = 4'h0;
    SS13[7][45] = 4'h0;
    SS13[8][45] = 4'h0;
    SS13[9][45] = 4'h0;
    SS13[10][45] = 4'h0;
    SS13[11][45] = 4'h0;
    SS13[12][45] = 4'h0;
    SS13[13][45] = 4'h0;
    SS13[14][45] = 4'h0;
    SS13[15][45] = 4'h0;
    SS13[16][45] = 4'h0;
    SS13[17][45] = 4'hC;
    SS13[18][45] = 4'hC;
    SS13[19][45] = 4'hC;
    SS13[20][45] = 4'hD;
    SS13[21][45] = 4'hD;
    SS13[22][45] = 4'hD;
    SS13[23][45] = 4'h0;
    SS13[24][45] = 4'h0;
    SS13[25][45] = 4'h0;
    SS13[26][45] = 4'h0;
    SS13[27][45] = 4'h0;
    SS13[28][45] = 4'h0;
    SS13[29][45] = 4'h0;
    SS13[30][45] = 4'h0;
    SS13[31][45] = 4'h0;
    SS13[32][45] = 4'h0;
    SS13[33][45] = 4'h0;
    SS13[34][45] = 4'h0;
    SS13[35][45] = 4'h0;
    SS13[36][45] = 4'h0;
    SS13[37][45] = 4'h0;
    SS13[38][45] = 4'h0;
    SS13[39][45] = 4'h0;
    SS13[40][45] = 4'h0;
    SS13[41][45] = 4'h0;
    SS13[42][45] = 4'h0;
    SS13[43][45] = 4'h0;
    SS13[44][45] = 4'h0;
    SS13[45][45] = 4'h0;
    SS13[46][45] = 4'h0;
    SS13[47][45] = 4'h0;
    SS13[0][46] = 4'h0;
    SS13[1][46] = 4'h0;
    SS13[2][46] = 4'h0;
    SS13[3][46] = 4'h0;
    SS13[4][46] = 4'h0;
    SS13[5][46] = 4'h0;
    SS13[6][46] = 4'h0;
    SS13[7][46] = 4'h0;
    SS13[8][46] = 4'h0;
    SS13[9][46] = 4'h0;
    SS13[10][46] = 4'h0;
    SS13[11][46] = 4'h0;
    SS13[12][46] = 4'h0;
    SS13[13][46] = 4'h0;
    SS13[14][46] = 4'h0;
    SS13[15][46] = 4'h0;
    SS13[16][46] = 4'h0;
    SS13[17][46] = 4'hC;
    SS13[18][46] = 4'hC;
    SS13[19][46] = 4'hC;
    SS13[20][46] = 4'hD;
    SS13[21][46] = 4'hD;
    SS13[22][46] = 4'hD;
    SS13[23][46] = 4'hD;
    SS13[24][46] = 4'h0;
    SS13[25][46] = 4'h0;
    SS13[26][46] = 4'h0;
    SS13[27][46] = 4'h0;
    SS13[28][46] = 4'h0;
    SS13[29][46] = 4'h0;
    SS13[30][46] = 4'h0;
    SS13[31][46] = 4'h0;
    SS13[32][46] = 4'h0;
    SS13[33][46] = 4'h0;
    SS13[34][46] = 4'h0;
    SS13[35][46] = 4'h0;
    SS13[36][46] = 4'h0;
    SS13[37][46] = 4'h0;
    SS13[38][46] = 4'h0;
    SS13[39][46] = 4'h0;
    SS13[40][46] = 4'h0;
    SS13[41][46] = 4'h0;
    SS13[42][46] = 4'h0;
    SS13[43][46] = 4'h0;
    SS13[44][46] = 4'h0;
    SS13[45][46] = 4'h0;
    SS13[46][46] = 4'h0;
    SS13[47][46] = 4'h0;
    SS13[0][47] = 4'h0;
    SS13[1][47] = 4'h0;
    SS13[2][47] = 4'h0;
    SS13[3][47] = 4'h0;
    SS13[4][47] = 4'h0;
    SS13[5][47] = 4'h0;
    SS13[6][47] = 4'h0;
    SS13[7][47] = 4'h0;
    SS13[8][47] = 4'h0;
    SS13[9][47] = 4'h0;
    SS13[10][47] = 4'h0;
    SS13[11][47] = 4'h0;
    SS13[12][47] = 4'h0;
    SS13[13][47] = 4'h0;
    SS13[14][47] = 4'h0;
    SS13[15][47] = 4'h0;
    SS13[16][47] = 4'h0;
    SS13[17][47] = 4'h0;
    SS13[18][47] = 4'hC;
    SS13[19][47] = 4'hC;
    SS13[20][47] = 4'hC;
    SS13[21][47] = 4'h0;
    SS13[22][47] = 4'h0;
    SS13[23][47] = 4'h0;
    SS13[24][47] = 4'h0;
    SS13[25][47] = 4'h0;
    SS13[26][47] = 4'h0;
    SS13[27][47] = 4'h0;
    SS13[28][47] = 4'h0;
    SS13[29][47] = 4'h0;
    SS13[30][47] = 4'h0;
    SS13[31][47] = 4'h0;
    SS13[32][47] = 4'h0;
    SS13[33][47] = 4'h0;
    SS13[34][47] = 4'h0;
    SS13[35][47] = 4'h0;
    SS13[36][47] = 4'h0;
    SS13[37][47] = 4'h0;
    SS13[38][47] = 4'h0;
    SS13[39][47] = 4'h0;
    SS13[40][47] = 4'h0;
    SS13[41][47] = 4'h0;
    SS13[42][47] = 4'h0;
    SS13[43][47] = 4'h0;
    SS13[44][47] = 4'h0;
    SS13[45][47] = 4'h0;
    SS13[46][47] = 4'h0;
    SS13[47][47] = 4'h0;
 
//SS 14
    SS14[0][0] = 4'h0;
    SS14[1][0] = 4'h0;
    SS14[2][0] = 4'h0;
    SS14[3][0] = 4'h0;
    SS14[4][0] = 4'h0;
    SS14[5][0] = 4'h0;
    SS14[6][0] = 4'h0;
    SS14[7][0] = 4'h0;
    SS14[8][0] = 4'h0;
    SS14[9][0] = 4'h0;
    SS14[10][0] = 4'h0;
    SS14[11][0] = 4'h0;
    SS14[12][0] = 4'h0;
    SS14[13][0] = 4'h0;
    SS14[14][0] = 4'h0;
    SS14[15][0] = 4'h0;
    SS14[16][0] = 4'h0;
    SS14[17][0] = 4'h0;
    SS14[18][0] = 4'h0;
    SS14[19][0] = 4'h0;
    SS14[20][0] = 4'h0;
    SS14[21][0] = 4'hC;
    SS14[22][0] = 4'hC;
    SS14[23][0] = 4'hC;
    SS14[24][0] = 4'hC;
    SS14[25][0] = 4'hC;
    SS14[26][0] = 4'hC;
    SS14[27][0] = 4'h0;
    SS14[28][0] = 4'h0;
    SS14[29][0] = 4'h0;
    SS14[30][0] = 4'h0;
    SS14[31][0] = 4'h0;
    SS14[32][0] = 4'h0;
    SS14[33][0] = 4'h0;
    SS14[34][0] = 4'h0;
    SS14[35][0] = 4'h0;
    SS14[36][0] = 4'h0;
    SS14[37][0] = 4'h0;
    SS14[38][0] = 4'h0;
    SS14[39][0] = 4'h0;
    SS14[40][0] = 4'h0;
    SS14[41][0] = 4'h0;
    SS14[42][0] = 4'h0;
    SS14[43][0] = 4'h0;
    SS14[44][0] = 4'h0;
    SS14[45][0] = 4'h0;
    SS14[46][0] = 4'h0;
    SS14[47][0] = 4'h0;
    SS14[0][1] = 4'h0;
    SS14[1][1] = 4'h0;
    SS14[2][1] = 4'h0;
    SS14[3][1] = 4'h0;
    SS14[4][1] = 4'h0;
    SS14[5][1] = 4'h0;
    SS14[6][1] = 4'h0;
    SS14[7][1] = 4'h0;
    SS14[8][1] = 4'h0;
    SS14[9][1] = 4'h0;
    SS14[10][1] = 4'h0;
    SS14[11][1] = 4'h0;
    SS14[12][1] = 4'h0;
    SS14[13][1] = 4'h0;
    SS14[14][1] = 4'h0;
    SS14[15][1] = 4'h0;
    SS14[16][1] = 4'h0;
    SS14[17][1] = 4'h0;
    SS14[18][1] = 4'h0;
    SS14[19][1] = 4'h0;
    SS14[20][1] = 4'h0;
    SS14[21][1] = 4'hC;
    SS14[22][1] = 4'hC;
    SS14[23][1] = 4'hC;
    SS14[24][1] = 4'hC;
    SS14[25][1] = 4'hC;
    SS14[26][1] = 4'hC;
    SS14[27][1] = 4'h0;
    SS14[28][1] = 4'h0;
    SS14[29][1] = 4'h0;
    SS14[30][1] = 4'h0;
    SS14[31][1] = 4'h0;
    SS14[32][1] = 4'h0;
    SS14[33][1] = 4'h0;
    SS14[34][1] = 4'h0;
    SS14[35][1] = 4'h0;
    SS14[36][1] = 4'h0;
    SS14[37][1] = 4'h0;
    SS14[38][1] = 4'h0;
    SS14[39][1] = 4'h0;
    SS14[40][1] = 4'h0;
    SS14[41][1] = 4'h0;
    SS14[42][1] = 4'h0;
    SS14[43][1] = 4'h0;
    SS14[44][1] = 4'h0;
    SS14[45][1] = 4'h0;
    SS14[46][1] = 4'h0;
    SS14[47][1] = 4'h0;
    SS14[0][2] = 4'h0;
    SS14[1][2] = 4'h0;
    SS14[2][2] = 4'h0;
    SS14[3][2] = 4'h0;
    SS14[4][2] = 4'h0;
    SS14[5][2] = 4'h0;
    SS14[6][2] = 4'h0;
    SS14[7][2] = 4'h0;
    SS14[8][2] = 4'h0;
    SS14[9][2] = 4'h0;
    SS14[10][2] = 4'h0;
    SS14[11][2] = 4'h0;
    SS14[12][2] = 4'h0;
    SS14[13][2] = 4'h0;
    SS14[14][2] = 4'h0;
    SS14[15][2] = 4'h0;
    SS14[16][2] = 4'h0;
    SS14[17][2] = 4'h0;
    SS14[18][2] = 4'h0;
    SS14[19][2] = 4'h0;
    SS14[20][2] = 4'h0;
    SS14[21][2] = 4'hC;
    SS14[22][2] = 4'hC;
    SS14[23][2] = 4'hC;
    SS14[24][2] = 4'hC;
    SS14[25][2] = 4'hC;
    SS14[26][2] = 4'hC;
    SS14[27][2] = 4'h0;
    SS14[28][2] = 4'h0;
    SS14[29][2] = 4'h0;
    SS14[30][2] = 4'h0;
    SS14[31][2] = 4'h0;
    SS14[32][2] = 4'h0;
    SS14[33][2] = 4'h0;
    SS14[34][2] = 4'h0;
    SS14[35][2] = 4'h0;
    SS14[36][2] = 4'h0;
    SS14[37][2] = 4'h0;
    SS14[38][2] = 4'h0;
    SS14[39][2] = 4'h0;
    SS14[40][2] = 4'h0;
    SS14[41][2] = 4'h0;
    SS14[42][2] = 4'h0;
    SS14[43][2] = 4'h0;
    SS14[44][2] = 4'h0;
    SS14[45][2] = 4'h0;
    SS14[46][2] = 4'h0;
    SS14[47][2] = 4'h0;
    SS14[0][3] = 4'h0;
    SS14[1][3] = 4'h0;
    SS14[2][3] = 4'h0;
    SS14[3][3] = 4'h0;
    SS14[4][3] = 4'h0;
    SS14[5][3] = 4'h0;
    SS14[6][3] = 4'h0;
    SS14[7][3] = 4'h0;
    SS14[8][3] = 4'h0;
    SS14[9][3] = 4'h0;
    SS14[10][3] = 4'h0;
    SS14[11][3] = 4'h0;
    SS14[12][3] = 4'h0;
    SS14[13][3] = 4'h0;
    SS14[14][3] = 4'h0;
    SS14[15][3] = 4'h0;
    SS14[16][3] = 4'h0;
    SS14[17][3] = 4'h0;
    SS14[18][3] = 4'h0;
    SS14[19][3] = 4'h0;
    SS14[20][3] = 4'h0;
    SS14[21][3] = 4'hC;
    SS14[22][3] = 4'hC;
    SS14[23][3] = 4'hC;
    SS14[24][3] = 4'hC;
    SS14[25][3] = 4'hC;
    SS14[26][3] = 4'hC;
    SS14[27][3] = 4'h0;
    SS14[28][3] = 4'h0;
    SS14[29][3] = 4'h0;
    SS14[30][3] = 4'h0;
    SS14[31][3] = 4'h0;
    SS14[32][3] = 4'h0;
    SS14[33][3] = 4'h0;
    SS14[34][3] = 4'h0;
    SS14[35][3] = 4'h0;
    SS14[36][3] = 4'h0;
    SS14[37][3] = 4'h0;
    SS14[38][3] = 4'h0;
    SS14[39][3] = 4'h0;
    SS14[40][3] = 4'h0;
    SS14[41][3] = 4'h0;
    SS14[42][3] = 4'h0;
    SS14[43][3] = 4'h0;
    SS14[44][3] = 4'h0;
    SS14[45][3] = 4'h0;
    SS14[46][3] = 4'h0;
    SS14[47][3] = 4'h0;
    SS14[0][4] = 4'h0;
    SS14[1][4] = 4'h0;
    SS14[2][4] = 4'h0;
    SS14[3][4] = 4'h0;
    SS14[4][4] = 4'h0;
    SS14[5][4] = 4'h0;
    SS14[6][4] = 4'h0;
    SS14[7][4] = 4'h0;
    SS14[8][4] = 4'h0;
    SS14[9][4] = 4'h0;
    SS14[10][4] = 4'h0;
    SS14[11][4] = 4'h0;
    SS14[12][4] = 4'h0;
    SS14[13][4] = 4'h0;
    SS14[14][4] = 4'h0;
    SS14[15][4] = 4'h0;
    SS14[16][4] = 4'h0;
    SS14[17][4] = 4'h0;
    SS14[18][4] = 4'h0;
    SS14[19][4] = 4'h0;
    SS14[20][4] = 4'h0;
    SS14[21][4] = 4'hC;
    SS14[22][4] = 4'hC;
    SS14[23][4] = 4'hC;
    SS14[24][4] = 4'hC;
    SS14[25][4] = 4'hC;
    SS14[26][4] = 4'hC;
    SS14[27][4] = 4'h0;
    SS14[28][4] = 4'h0;
    SS14[29][4] = 4'h0;
    SS14[30][4] = 4'h0;
    SS14[31][4] = 4'h0;
    SS14[32][4] = 4'h0;
    SS14[33][4] = 4'h0;
    SS14[34][4] = 4'h0;
    SS14[35][4] = 4'h0;
    SS14[36][4] = 4'h0;
    SS14[37][4] = 4'h0;
    SS14[38][4] = 4'h0;
    SS14[39][4] = 4'h0;
    SS14[40][4] = 4'h0;
    SS14[41][4] = 4'h0;
    SS14[42][4] = 4'h0;
    SS14[43][4] = 4'h0;
    SS14[44][4] = 4'h0;
    SS14[45][4] = 4'h0;
    SS14[46][4] = 4'h0;
    SS14[47][4] = 4'h0;
    SS14[0][5] = 4'h0;
    SS14[1][5] = 4'h0;
    SS14[2][5] = 4'h0;
    SS14[3][5] = 4'h0;
    SS14[4][5] = 4'h0;
    SS14[5][5] = 4'h0;
    SS14[6][5] = 4'h0;
    SS14[7][5] = 4'h0;
    SS14[8][5] = 4'h0;
    SS14[9][5] = 4'h0;
    SS14[10][5] = 4'h0;
    SS14[11][5] = 4'h0;
    SS14[12][5] = 4'h0;
    SS14[13][5] = 4'h0;
    SS14[14][5] = 4'h0;
    SS14[15][5] = 4'h0;
    SS14[16][5] = 4'h0;
    SS14[17][5] = 4'h0;
    SS14[18][5] = 4'h0;
    SS14[19][5] = 4'h0;
    SS14[20][5] = 4'h0;
    SS14[21][5] = 4'hC;
    SS14[22][5] = 4'hC;
    SS14[23][5] = 4'hC;
    SS14[24][5] = 4'hC;
    SS14[25][5] = 4'hC;
    SS14[26][5] = 4'hC;
    SS14[27][5] = 4'h0;
    SS14[28][5] = 4'h0;
    SS14[29][5] = 4'h0;
    SS14[30][5] = 4'h0;
    SS14[31][5] = 4'h0;
    SS14[32][5] = 4'h0;
    SS14[33][5] = 4'h0;
    SS14[34][5] = 4'h0;
    SS14[35][5] = 4'h0;
    SS14[36][5] = 4'h0;
    SS14[37][5] = 4'h0;
    SS14[38][5] = 4'h0;
    SS14[39][5] = 4'h0;
    SS14[40][5] = 4'h0;
    SS14[41][5] = 4'h0;
    SS14[42][5] = 4'h0;
    SS14[43][5] = 4'h0;
    SS14[44][5] = 4'h0;
    SS14[45][5] = 4'h0;
    SS14[46][5] = 4'h0;
    SS14[47][5] = 4'h0;
    SS14[0][6] = 4'h0;
    SS14[1][6] = 4'h0;
    SS14[2][6] = 4'h0;
    SS14[3][6] = 4'h0;
    SS14[4][6] = 4'h0;
    SS14[5][6] = 4'h0;
    SS14[6][6] = 4'h0;
    SS14[7][6] = 4'h0;
    SS14[8][6] = 4'h0;
    SS14[9][6] = 4'h0;
    SS14[10][6] = 4'h0;
    SS14[11][6] = 4'h0;
    SS14[12][6] = 4'h0;
    SS14[13][6] = 4'h0;
    SS14[14][6] = 4'h0;
    SS14[15][6] = 4'h0;
    SS14[16][6] = 4'h0;
    SS14[17][6] = 4'h0;
    SS14[18][6] = 4'hD;
    SS14[19][6] = 4'hD;
    SS14[20][6] = 4'hD;
    SS14[21][6] = 4'hC;
    SS14[22][6] = 4'hC;
    SS14[23][6] = 4'hC;
    SS14[24][6] = 4'hC;
    SS14[25][6] = 4'hC;
    SS14[26][6] = 4'hC;
    SS14[27][6] = 4'hD;
    SS14[28][6] = 4'hD;
    SS14[29][6] = 4'hD;
    SS14[30][6] = 4'h0;
    SS14[31][6] = 4'h0;
    SS14[32][6] = 4'h0;
    SS14[33][6] = 4'h0;
    SS14[34][6] = 4'h0;
    SS14[35][6] = 4'h0;
    SS14[36][6] = 4'h0;
    SS14[37][6] = 4'h0;
    SS14[38][6] = 4'h0;
    SS14[39][6] = 4'h0;
    SS14[40][6] = 4'h0;
    SS14[41][6] = 4'h0;
    SS14[42][6] = 4'h0;
    SS14[43][6] = 4'h0;
    SS14[44][6] = 4'h0;
    SS14[45][6] = 4'h0;
    SS14[46][6] = 4'h0;
    SS14[47][6] = 4'h0;
    SS14[0][7] = 4'h0;
    SS14[1][7] = 4'h0;
    SS14[2][7] = 4'h0;
    SS14[3][7] = 4'h0;
    SS14[4][7] = 4'h0;
    SS14[5][7] = 4'h0;
    SS14[6][7] = 4'h0;
    SS14[7][7] = 4'h0;
    SS14[8][7] = 4'h0;
    SS14[9][7] = 4'h0;
    SS14[10][7] = 4'h0;
    SS14[11][7] = 4'h0;
    SS14[12][7] = 4'h0;
    SS14[13][7] = 4'h0;
    SS14[14][7] = 4'h0;
    SS14[15][7] = 4'h0;
    SS14[16][7] = 4'h0;
    SS14[17][7] = 4'h0;
    SS14[18][7] = 4'hD;
    SS14[19][7] = 4'hD;
    SS14[20][7] = 4'hD;
    SS14[21][7] = 4'hC;
    SS14[22][7] = 4'hC;
    SS14[23][7] = 4'hC;
    SS14[24][7] = 4'hC;
    SS14[25][7] = 4'hC;
    SS14[26][7] = 4'hC;
    SS14[27][7] = 4'hD;
    SS14[28][7] = 4'hD;
    SS14[29][7] = 4'hD;
    SS14[30][7] = 4'h0;
    SS14[31][7] = 4'h0;
    SS14[32][7] = 4'h0;
    SS14[33][7] = 4'h0;
    SS14[34][7] = 4'h0;
    SS14[35][7] = 4'h0;
    SS14[36][7] = 4'h0;
    SS14[37][7] = 4'h0;
    SS14[38][7] = 4'h0;
    SS14[39][7] = 4'h0;
    SS14[40][7] = 4'h0;
    SS14[41][7] = 4'h0;
    SS14[42][7] = 4'h0;
    SS14[43][7] = 4'h0;
    SS14[44][7] = 4'h0;
    SS14[45][7] = 4'h0;
    SS14[46][7] = 4'h0;
    SS14[47][7] = 4'h0;
    SS14[0][8] = 4'h0;
    SS14[1][8] = 4'h0;
    SS14[2][8] = 4'h0;
    SS14[3][8] = 4'h0;
    SS14[4][8] = 4'h0;
    SS14[5][8] = 4'h0;
    SS14[6][8] = 4'h0;
    SS14[7][8] = 4'h0;
    SS14[8][8] = 4'h0;
    SS14[9][8] = 4'h0;
    SS14[10][8] = 4'h0;
    SS14[11][8] = 4'h0;
    SS14[12][8] = 4'h0;
    SS14[13][8] = 4'h0;
    SS14[14][8] = 4'h0;
    SS14[15][8] = 4'h0;
    SS14[16][8] = 4'h0;
    SS14[17][8] = 4'h0;
    SS14[18][8] = 4'hD;
    SS14[19][8] = 4'hD;
    SS14[20][8] = 4'hD;
    SS14[21][8] = 4'hC;
    SS14[22][8] = 4'hC;
    SS14[23][8] = 4'hC;
    SS14[24][8] = 4'hC;
    SS14[25][8] = 4'hC;
    SS14[26][8] = 4'hC;
    SS14[27][8] = 4'hD;
    SS14[28][8] = 4'hD;
    SS14[29][8] = 4'hD;
    SS14[30][8] = 4'h0;
    SS14[31][8] = 4'h0;
    SS14[32][8] = 4'h0;
    SS14[33][8] = 4'h0;
    SS14[34][8] = 4'h0;
    SS14[35][8] = 4'h0;
    SS14[36][8] = 4'h0;
    SS14[37][8] = 4'h0;
    SS14[38][8] = 4'h0;
    SS14[39][8] = 4'h0;
    SS14[40][8] = 4'h0;
    SS14[41][8] = 4'h0;
    SS14[42][8] = 4'h0;
    SS14[43][8] = 4'h0;
    SS14[44][8] = 4'h0;
    SS14[45][8] = 4'h0;
    SS14[46][8] = 4'h0;
    SS14[47][8] = 4'h0;
    SS14[0][9] = 4'h0;
    SS14[1][9] = 4'h0;
    SS14[2][9] = 4'h0;
    SS14[3][9] = 4'h0;
    SS14[4][9] = 4'h0;
    SS14[5][9] = 4'h0;
    SS14[6][9] = 4'h0;
    SS14[7][9] = 4'h0;
    SS14[8][9] = 4'h0;
    SS14[9][9] = 4'h0;
    SS14[10][9] = 4'h0;
    SS14[11][9] = 4'h0;
    SS14[12][9] = 4'h0;
    SS14[13][9] = 4'h0;
    SS14[14][9] = 4'h0;
    SS14[15][9] = 4'h0;
    SS14[16][9] = 4'h0;
    SS14[17][9] = 4'h0;
    SS14[18][9] = 4'hD;
    SS14[19][9] = 4'hD;
    SS14[20][9] = 4'hD;
    SS14[21][9] = 4'hC;
    SS14[22][9] = 4'hC;
    SS14[23][9] = 4'hC;
    SS14[24][9] = 4'hC;
    SS14[25][9] = 4'hC;
    SS14[26][9] = 4'hC;
    SS14[27][9] = 4'hD;
    SS14[28][9] = 4'hD;
    SS14[29][9] = 4'hD;
    SS14[30][9] = 4'h0;
    SS14[31][9] = 4'h0;
    SS14[32][9] = 4'h0;
    SS14[33][9] = 4'h0;
    SS14[34][9] = 4'h0;
    SS14[35][9] = 4'h0;
    SS14[36][9] = 4'h0;
    SS14[37][9] = 4'h0;
    SS14[38][9] = 4'h0;
    SS14[39][9] = 4'h0;
    SS14[40][9] = 4'h0;
    SS14[41][9] = 4'h0;
    SS14[42][9] = 4'h0;
    SS14[43][9] = 4'h0;
    SS14[44][9] = 4'h0;
    SS14[45][9] = 4'h0;
    SS14[46][9] = 4'h0;
    SS14[47][9] = 4'h0;
    SS14[0][10] = 4'h0;
    SS14[1][10] = 4'h0;
    SS14[2][10] = 4'h0;
    SS14[3][10] = 4'h0;
    SS14[4][10] = 4'h0;
    SS14[5][10] = 4'h0;
    SS14[6][10] = 4'h0;
    SS14[7][10] = 4'h0;
    SS14[8][10] = 4'h0;
    SS14[9][10] = 4'h0;
    SS14[10][10] = 4'h0;
    SS14[11][10] = 4'h0;
    SS14[12][10] = 4'h0;
    SS14[13][10] = 4'h0;
    SS14[14][10] = 4'h0;
    SS14[15][10] = 4'h0;
    SS14[16][10] = 4'h0;
    SS14[17][10] = 4'h0;
    SS14[18][10] = 4'hD;
    SS14[19][10] = 4'hD;
    SS14[20][10] = 4'hD;
    SS14[21][10] = 4'hC;
    SS14[22][10] = 4'hC;
    SS14[23][10] = 4'hC;
    SS14[24][10] = 4'hC;
    SS14[25][10] = 4'hC;
    SS14[26][10] = 4'hC;
    SS14[27][10] = 4'hD;
    SS14[28][10] = 4'hD;
    SS14[29][10] = 4'hD;
    SS14[30][10] = 4'h0;
    SS14[31][10] = 4'h0;
    SS14[32][10] = 4'h0;
    SS14[33][10] = 4'h0;
    SS14[34][10] = 4'h0;
    SS14[35][10] = 4'h0;
    SS14[36][10] = 4'h0;
    SS14[37][10] = 4'h0;
    SS14[38][10] = 4'h0;
    SS14[39][10] = 4'h0;
    SS14[40][10] = 4'h0;
    SS14[41][10] = 4'h0;
    SS14[42][10] = 4'h0;
    SS14[43][10] = 4'h0;
    SS14[44][10] = 4'h0;
    SS14[45][10] = 4'h0;
    SS14[46][10] = 4'h0;
    SS14[47][10] = 4'h0;
    SS14[0][11] = 4'h0;
    SS14[1][11] = 4'h0;
    SS14[2][11] = 4'h0;
    SS14[3][11] = 4'h0;
    SS14[4][11] = 4'h0;
    SS14[5][11] = 4'h0;
    SS14[6][11] = 4'h0;
    SS14[7][11] = 4'h0;
    SS14[8][11] = 4'h0;
    SS14[9][11] = 4'h0;
    SS14[10][11] = 4'h0;
    SS14[11][11] = 4'h0;
    SS14[12][11] = 4'h0;
    SS14[13][11] = 4'h0;
    SS14[14][11] = 4'h0;
    SS14[15][11] = 4'h0;
    SS14[16][11] = 4'h0;
    SS14[17][11] = 4'h0;
    SS14[18][11] = 4'hD;
    SS14[19][11] = 4'hD;
    SS14[20][11] = 4'hD;
    SS14[21][11] = 4'hC;
    SS14[22][11] = 4'hC;
    SS14[23][11] = 4'hC;
    SS14[24][11] = 4'hC;
    SS14[25][11] = 4'hC;
    SS14[26][11] = 4'hC;
    SS14[27][11] = 4'hD;
    SS14[28][11] = 4'hD;
    SS14[29][11] = 4'hD;
    SS14[30][11] = 4'h0;
    SS14[31][11] = 4'h0;
    SS14[32][11] = 4'h0;
    SS14[33][11] = 4'h0;
    SS14[34][11] = 4'h0;
    SS14[35][11] = 4'h0;
    SS14[36][11] = 4'h0;
    SS14[37][11] = 4'h0;
    SS14[38][11] = 4'h0;
    SS14[39][11] = 4'h0;
    SS14[40][11] = 4'h0;
    SS14[41][11] = 4'h0;
    SS14[42][11] = 4'h0;
    SS14[43][11] = 4'h0;
    SS14[44][11] = 4'h0;
    SS14[45][11] = 4'h0;
    SS14[46][11] = 4'h0;
    SS14[47][11] = 4'h0;
    SS14[0][12] = 4'h0;
    SS14[1][12] = 4'h0;
    SS14[2][12] = 4'h0;
    SS14[3][12] = 4'h0;
    SS14[4][12] = 4'h0;
    SS14[5][12] = 4'h0;
    SS14[6][12] = 4'h0;
    SS14[7][12] = 4'h0;
    SS14[8][12] = 4'h0;
    SS14[9][12] = 4'h0;
    SS14[10][12] = 4'h0;
    SS14[11][12] = 4'h0;
    SS14[12][12] = 4'h0;
    SS14[13][12] = 4'h0;
    SS14[14][12] = 4'h0;
    SS14[15][12] = 4'h0;
    SS14[16][12] = 4'h0;
    SS14[17][12] = 4'h0;
    SS14[18][12] = 4'hD;
    SS14[19][12] = 4'hD;
    SS14[20][12] = 4'hD;
    SS14[21][12] = 4'hC;
    SS14[22][12] = 4'hC;
    SS14[23][12] = 4'hC;
    SS14[24][12] = 4'hC;
    SS14[25][12] = 4'hC;
    SS14[26][12] = 4'hC;
    SS14[27][12] = 4'hD;
    SS14[28][12] = 4'hD;
    SS14[29][12] = 4'hD;
    SS14[30][12] = 4'h0;
    SS14[31][12] = 4'h0;
    SS14[32][12] = 4'h0;
    SS14[33][12] = 4'h0;
    SS14[34][12] = 4'h0;
    SS14[35][12] = 4'h0;
    SS14[36][12] = 4'h0;
    SS14[37][12] = 4'h0;
    SS14[38][12] = 4'h0;
    SS14[39][12] = 4'h0;
    SS14[40][12] = 4'h0;
    SS14[41][12] = 4'h0;
    SS14[42][12] = 4'h0;
    SS14[43][12] = 4'h0;
    SS14[44][12] = 4'h0;
    SS14[45][12] = 4'h0;
    SS14[46][12] = 4'h0;
    SS14[47][12] = 4'h0;
    SS14[0][13] = 4'h0;
    SS14[1][13] = 4'h0;
    SS14[2][13] = 4'h0;
    SS14[3][13] = 4'h0;
    SS14[4][13] = 4'h0;
    SS14[5][13] = 4'h0;
    SS14[6][13] = 4'h0;
    SS14[7][13] = 4'h0;
    SS14[8][13] = 4'h0;
    SS14[9][13] = 4'h0;
    SS14[10][13] = 4'h0;
    SS14[11][13] = 4'h0;
    SS14[12][13] = 4'h0;
    SS14[13][13] = 4'h0;
    SS14[14][13] = 4'h0;
    SS14[15][13] = 4'h0;
    SS14[16][13] = 4'h0;
    SS14[17][13] = 4'h0;
    SS14[18][13] = 4'hD;
    SS14[19][13] = 4'hD;
    SS14[20][13] = 4'hD;
    SS14[21][13] = 4'hC;
    SS14[22][13] = 4'hC;
    SS14[23][13] = 4'hC;
    SS14[24][13] = 4'hC;
    SS14[25][13] = 4'hC;
    SS14[26][13] = 4'hC;
    SS14[27][13] = 4'hD;
    SS14[28][13] = 4'hD;
    SS14[29][13] = 4'hD;
    SS14[30][13] = 4'h0;
    SS14[31][13] = 4'h0;
    SS14[32][13] = 4'h0;
    SS14[33][13] = 4'h0;
    SS14[34][13] = 4'h0;
    SS14[35][13] = 4'h0;
    SS14[36][13] = 4'h0;
    SS14[37][13] = 4'h0;
    SS14[38][13] = 4'h0;
    SS14[39][13] = 4'h0;
    SS14[40][13] = 4'h0;
    SS14[41][13] = 4'h0;
    SS14[42][13] = 4'h0;
    SS14[43][13] = 4'h0;
    SS14[44][13] = 4'h0;
    SS14[45][13] = 4'h0;
    SS14[46][13] = 4'h0;
    SS14[47][13] = 4'h0;
    SS14[0][14] = 4'h0;
    SS14[1][14] = 4'h0;
    SS14[2][14] = 4'h0;
    SS14[3][14] = 4'h0;
    SS14[4][14] = 4'h0;
    SS14[5][14] = 4'h0;
    SS14[6][14] = 4'h0;
    SS14[7][14] = 4'h0;
    SS14[8][14] = 4'h0;
    SS14[9][14] = 4'h0;
    SS14[10][14] = 4'h0;
    SS14[11][14] = 4'h0;
    SS14[12][14] = 4'h0;
    SS14[13][14] = 4'h0;
    SS14[14][14] = 4'h0;
    SS14[15][14] = 4'h0;
    SS14[16][14] = 4'h0;
    SS14[17][14] = 4'h0;
    SS14[18][14] = 4'hD;
    SS14[19][14] = 4'hD;
    SS14[20][14] = 4'hD;
    SS14[21][14] = 4'hC;
    SS14[22][14] = 4'hC;
    SS14[23][14] = 4'hC;
    SS14[24][14] = 4'hC;
    SS14[25][14] = 4'hC;
    SS14[26][14] = 4'hC;
    SS14[27][14] = 4'hD;
    SS14[28][14] = 4'hD;
    SS14[29][14] = 4'hD;
    SS14[30][14] = 4'h0;
    SS14[31][14] = 4'h0;
    SS14[32][14] = 4'h0;
    SS14[33][14] = 4'h0;
    SS14[34][14] = 4'h0;
    SS14[35][14] = 4'h0;
    SS14[36][14] = 4'h0;
    SS14[37][14] = 4'h0;
    SS14[38][14] = 4'h0;
    SS14[39][14] = 4'h0;
    SS14[40][14] = 4'h0;
    SS14[41][14] = 4'h0;
    SS14[42][14] = 4'h0;
    SS14[43][14] = 4'h0;
    SS14[44][14] = 4'h0;
    SS14[45][14] = 4'h0;
    SS14[46][14] = 4'h0;
    SS14[47][14] = 4'h0;
    SS14[0][15] = 4'h0;
    SS14[1][15] = 4'h0;
    SS14[2][15] = 4'h0;
    SS14[3][15] = 4'h0;
    SS14[4][15] = 4'h0;
    SS14[5][15] = 4'h0;
    SS14[6][15] = 4'h0;
    SS14[7][15] = 4'h0;
    SS14[8][15] = 4'h0;
    SS14[9][15] = 4'h0;
    SS14[10][15] = 4'h0;
    SS14[11][15] = 4'h0;
    SS14[12][15] = 4'h0;
    SS14[13][15] = 4'h0;
    SS14[14][15] = 4'h0;
    SS14[15][15] = 4'h0;
    SS14[16][15] = 4'h0;
    SS14[17][15] = 4'h0;
    SS14[18][15] = 4'hC;
    SS14[19][15] = 4'hC;
    SS14[20][15] = 4'hC;
    SS14[21][15] = 4'hC;
    SS14[22][15] = 4'hC;
    SS14[23][15] = 4'hC;
    SS14[24][15] = 4'hC;
    SS14[25][15] = 4'hC;
    SS14[26][15] = 4'hC;
    SS14[27][15] = 4'hC;
    SS14[28][15] = 4'hC;
    SS14[29][15] = 4'hC;
    SS14[30][15] = 4'h0;
    SS14[31][15] = 4'h0;
    SS14[32][15] = 4'h0;
    SS14[33][15] = 4'h0;
    SS14[34][15] = 4'h0;
    SS14[35][15] = 4'h0;
    SS14[36][15] = 4'h0;
    SS14[37][15] = 4'h0;
    SS14[38][15] = 4'h0;
    SS14[39][15] = 4'h0;
    SS14[40][15] = 4'h0;
    SS14[41][15] = 4'h0;
    SS14[42][15] = 4'h0;
    SS14[43][15] = 4'h0;
    SS14[44][15] = 4'h0;
    SS14[45][15] = 4'h0;
    SS14[46][15] = 4'h0;
    SS14[47][15] = 4'h0;
    SS14[0][16] = 4'h0;
    SS14[1][16] = 4'h0;
    SS14[2][16] = 4'h0;
    SS14[3][16] = 4'h0;
    SS14[4][16] = 4'h0;
    SS14[5][16] = 4'h0;
    SS14[6][16] = 4'h0;
    SS14[7][16] = 4'h0;
    SS14[8][16] = 4'h0;
    SS14[9][16] = 4'h0;
    SS14[10][16] = 4'h0;
    SS14[11][16] = 4'h0;
    SS14[12][16] = 4'h0;
    SS14[13][16] = 4'h0;
    SS14[14][16] = 4'h0;
    SS14[15][16] = 4'h0;
    SS14[16][16] = 4'h0;
    SS14[17][16] = 4'h0;
    SS14[18][16] = 4'hC;
    SS14[19][16] = 4'hC;
    SS14[20][16] = 4'hC;
    SS14[21][16] = 4'hC;
    SS14[22][16] = 4'hC;
    SS14[23][16] = 4'hC;
    SS14[24][16] = 4'hC;
    SS14[25][16] = 4'hC;
    SS14[26][16] = 4'hC;
    SS14[27][16] = 4'hC;
    SS14[28][16] = 4'hC;
    SS14[29][16] = 4'hC;
    SS14[30][16] = 4'h0;
    SS14[31][16] = 4'h0;
    SS14[32][16] = 4'h0;
    SS14[33][16] = 4'h0;
    SS14[34][16] = 4'h0;
    SS14[35][16] = 4'h0;
    SS14[36][16] = 4'h0;
    SS14[37][16] = 4'h0;
    SS14[38][16] = 4'h0;
    SS14[39][16] = 4'h0;
    SS14[40][16] = 4'h0;
    SS14[41][16] = 4'h0;
    SS14[42][16] = 4'h0;
    SS14[43][16] = 4'h0;
    SS14[44][16] = 4'h0;
    SS14[45][16] = 4'h0;
    SS14[46][16] = 4'h0;
    SS14[47][16] = 4'h0;
    SS14[0][17] = 4'h0;
    SS14[1][17] = 4'h0;
    SS14[2][17] = 4'h0;
    SS14[3][17] = 4'h0;
    SS14[4][17] = 4'h0;
    SS14[5][17] = 4'h0;
    SS14[6][17] = 4'h0;
    SS14[7][17] = 4'h0;
    SS14[8][17] = 4'h0;
    SS14[9][17] = 4'h0;
    SS14[10][17] = 4'h0;
    SS14[11][17] = 4'h0;
    SS14[12][17] = 4'h0;
    SS14[13][17] = 4'h0;
    SS14[14][17] = 4'h0;
    SS14[15][17] = 4'h0;
    SS14[16][17] = 4'h0;
    SS14[17][17] = 4'h0;
    SS14[18][17] = 4'hC;
    SS14[19][17] = 4'hC;
    SS14[20][17] = 4'hC;
    SS14[21][17] = 4'hC;
    SS14[22][17] = 4'hC;
    SS14[23][17] = 4'hC;
    SS14[24][17] = 4'hC;
    SS14[25][17] = 4'hC;
    SS14[26][17] = 4'hC;
    SS14[27][17] = 4'hC;
    SS14[28][17] = 4'hC;
    SS14[29][17] = 4'hC;
    SS14[30][17] = 4'h0;
    SS14[31][17] = 4'h0;
    SS14[32][17] = 4'h0;
    SS14[33][17] = 4'h0;
    SS14[34][17] = 4'h0;
    SS14[35][17] = 4'h0;
    SS14[36][17] = 4'h0;
    SS14[37][17] = 4'h0;
    SS14[38][17] = 4'h0;
    SS14[39][17] = 4'h0;
    SS14[40][17] = 4'h0;
    SS14[41][17] = 4'h0;
    SS14[42][17] = 4'h0;
    SS14[43][17] = 4'h0;
    SS14[44][17] = 4'h0;
    SS14[45][17] = 4'h0;
    SS14[46][17] = 4'h0;
    SS14[47][17] = 4'h0;
    SS14[0][18] = 4'h0;
    SS14[1][18] = 4'h0;
    SS14[2][18] = 4'h0;
    SS14[3][18] = 4'h0;
    SS14[4][18] = 4'h0;
    SS14[5][18] = 4'h0;
    SS14[6][18] = 4'h0;
    SS14[7][18] = 4'h0;
    SS14[8][18] = 4'h0;
    SS14[9][18] = 4'h0;
    SS14[10][18] = 4'h0;
    SS14[11][18] = 4'h0;
    SS14[12][18] = 4'h3;
    SS14[13][18] = 4'h3;
    SS14[14][18] = 4'h3;
    SS14[15][18] = 4'hD;
    SS14[16][18] = 4'hD;
    SS14[17][18] = 4'hD;
    SS14[18][18] = 4'hD;
    SS14[19][18] = 4'hD;
    SS14[20][18] = 4'hD;
    SS14[21][18] = 4'hA;
    SS14[22][18] = 4'hA;
    SS14[23][18] = 4'hA;
    SS14[24][18] = 4'hA;
    SS14[25][18] = 4'hA;
    SS14[26][18] = 4'hA;
    SS14[27][18] = 4'hD;
    SS14[28][18] = 4'hD;
    SS14[29][18] = 4'hD;
    SS14[30][18] = 4'hD;
    SS14[31][18] = 4'hD;
    SS14[32][18] = 4'hD;
    SS14[33][18] = 4'h3;
    SS14[34][18] = 4'h3;
    SS14[35][18] = 4'h3;
    SS14[36][18] = 4'h0;
    SS14[37][18] = 4'h0;
    SS14[38][18] = 4'h0;
    SS14[39][18] = 4'h0;
    SS14[40][18] = 4'h0;
    SS14[41][18] = 4'h0;
    SS14[42][18] = 4'h0;
    SS14[43][18] = 4'h0;
    SS14[44][18] = 4'h0;
    SS14[45][18] = 4'h0;
    SS14[46][18] = 4'h0;
    SS14[47][18] = 4'h0;
    SS14[0][19] = 4'h0;
    SS14[1][19] = 4'h0;
    SS14[2][19] = 4'h0;
    SS14[3][19] = 4'h0;
    SS14[4][19] = 4'h0;
    SS14[5][19] = 4'h0;
    SS14[6][19] = 4'h0;
    SS14[7][19] = 4'h0;
    SS14[8][19] = 4'h0;
    SS14[9][19] = 4'h0;
    SS14[10][19] = 4'h0;
    SS14[11][19] = 4'h0;
    SS14[12][19] = 4'h3;
    SS14[13][19] = 4'h3;
    SS14[14][19] = 4'h3;
    SS14[15][19] = 4'hD;
    SS14[16][19] = 4'hD;
    SS14[17][19] = 4'hD;
    SS14[18][19] = 4'hD;
    SS14[19][19] = 4'hD;
    SS14[20][19] = 4'hD;
    SS14[21][19] = 4'hA;
    SS14[22][19] = 4'hA;
    SS14[23][19] = 4'hA;
    SS14[24][19] = 4'hA;
    SS14[25][19] = 4'hA;
    SS14[26][19] = 4'hA;
    SS14[27][19] = 4'hD;
    SS14[28][19] = 4'hD;
    SS14[29][19] = 4'hD;
    SS14[30][19] = 4'hD;
    SS14[31][19] = 4'hD;
    SS14[32][19] = 4'hD;
    SS14[33][19] = 4'h3;
    SS14[34][19] = 4'h3;
    SS14[35][19] = 4'h3;
    SS14[36][19] = 4'h0;
    SS14[37][19] = 4'h0;
    SS14[38][19] = 4'h0;
    SS14[39][19] = 4'h0;
    SS14[40][19] = 4'h0;
    SS14[41][19] = 4'h0;
    SS14[42][19] = 4'h0;
    SS14[43][19] = 4'h0;
    SS14[44][19] = 4'h0;
    SS14[45][19] = 4'h0;
    SS14[46][19] = 4'h0;
    SS14[47][19] = 4'h0;
    SS14[0][20] = 4'h0;
    SS14[1][20] = 4'h0;
    SS14[2][20] = 4'h0;
    SS14[3][20] = 4'h0;
    SS14[4][20] = 4'h0;
    SS14[5][20] = 4'h0;
    SS14[6][20] = 4'h0;
    SS14[7][20] = 4'h0;
    SS14[8][20] = 4'h0;
    SS14[9][20] = 4'h0;
    SS14[10][20] = 4'h0;
    SS14[11][20] = 4'h0;
    SS14[12][20] = 4'h3;
    SS14[13][20] = 4'h3;
    SS14[14][20] = 4'h3;
    SS14[15][20] = 4'hD;
    SS14[16][20] = 4'hD;
    SS14[17][20] = 4'hD;
    SS14[18][20] = 4'hD;
    SS14[19][20] = 4'hD;
    SS14[20][20] = 4'hD;
    SS14[21][20] = 4'hA;
    SS14[22][20] = 4'hA;
    SS14[23][20] = 4'hA;
    SS14[24][20] = 4'hA;
    SS14[25][20] = 4'hA;
    SS14[26][20] = 4'hA;
    SS14[27][20] = 4'hD;
    SS14[28][20] = 4'hD;
    SS14[29][20] = 4'hD;
    SS14[30][20] = 4'hD;
    SS14[31][20] = 4'hD;
    SS14[32][20] = 4'hD;
    SS14[33][20] = 4'h3;
    SS14[34][20] = 4'h3;
    SS14[35][20] = 4'h3;
    SS14[36][20] = 4'h0;
    SS14[37][20] = 4'h0;
    SS14[38][20] = 4'h0;
    SS14[39][20] = 4'h0;
    SS14[40][20] = 4'h0;
    SS14[41][20] = 4'h0;
    SS14[42][20] = 4'h0;
    SS14[43][20] = 4'h0;
    SS14[44][20] = 4'h0;
    SS14[45][20] = 4'h0;
    SS14[46][20] = 4'h0;
    SS14[47][20] = 4'h0;
    SS14[0][21] = 4'h0;
    SS14[1][21] = 4'h0;
    SS14[2][21] = 4'h0;
    SS14[3][21] = 4'h0;
    SS14[4][21] = 4'h0;
    SS14[5][21] = 4'h0;
    SS14[6][21] = 4'h0;
    SS14[7][21] = 4'h0;
    SS14[8][21] = 4'h0;
    SS14[9][21] = 4'h0;
    SS14[10][21] = 4'h0;
    SS14[11][21] = 4'h0;
    SS14[12][21] = 4'hD;
    SS14[13][21] = 4'hD;
    SS14[14][21] = 4'hD;
    SS14[15][21] = 4'hD;
    SS14[16][21] = 4'hD;
    SS14[17][21] = 4'hD;
    SS14[18][21] = 4'hC;
    SS14[19][21] = 4'hC;
    SS14[20][21] = 4'hC;
    SS14[21][21] = 4'hD;
    SS14[22][21] = 4'hD;
    SS14[23][21] = 4'hD;
    SS14[24][21] = 4'hD;
    SS14[25][21] = 4'hD;
    SS14[26][21] = 4'hD;
    SS14[27][21] = 4'hC;
    SS14[28][21] = 4'hC;
    SS14[29][21] = 4'hC;
    SS14[30][21] = 4'hD;
    SS14[31][21] = 4'hD;
    SS14[32][21] = 4'hD;
    SS14[33][21] = 4'hD;
    SS14[34][21] = 4'hD;
    SS14[35][21] = 4'hD;
    SS14[36][21] = 4'h0;
    SS14[37][21] = 4'h0;
    SS14[38][21] = 4'h0;
    SS14[39][21] = 4'h0;
    SS14[40][21] = 4'h0;
    SS14[41][21] = 4'h0;
    SS14[42][21] = 4'h0;
    SS14[43][21] = 4'h0;
    SS14[44][21] = 4'h0;
    SS14[45][21] = 4'h0;
    SS14[46][21] = 4'h0;
    SS14[47][21] = 4'h0;
    SS14[0][22] = 4'h0;
    SS14[1][22] = 4'h0;
    SS14[2][22] = 4'h0;
    SS14[3][22] = 4'h0;
    SS14[4][22] = 4'h0;
    SS14[5][22] = 4'h0;
    SS14[6][22] = 4'h0;
    SS14[7][22] = 4'h0;
    SS14[8][22] = 4'h0;
    SS14[9][22] = 4'h0;
    SS14[10][22] = 4'h0;
    SS14[11][22] = 4'h0;
    SS14[12][22] = 4'hD;
    SS14[13][22] = 4'hD;
    SS14[14][22] = 4'hD;
    SS14[15][22] = 4'hD;
    SS14[16][22] = 4'hD;
    SS14[17][22] = 4'hD;
    SS14[18][22] = 4'hC;
    SS14[19][22] = 4'hC;
    SS14[20][22] = 4'hC;
    SS14[21][22] = 4'hD;
    SS14[22][22] = 4'hD;
    SS14[23][22] = 4'hD;
    SS14[24][22] = 4'hD;
    SS14[25][22] = 4'hD;
    SS14[26][22] = 4'hD;
    SS14[27][22] = 4'hC;
    SS14[28][22] = 4'hC;
    SS14[29][22] = 4'hC;
    SS14[30][22] = 4'hD;
    SS14[31][22] = 4'hD;
    SS14[32][22] = 4'hD;
    SS14[33][22] = 4'hD;
    SS14[34][22] = 4'hD;
    SS14[35][22] = 4'hD;
    SS14[36][22] = 4'h0;
    SS14[37][22] = 4'h0;
    SS14[38][22] = 4'h0;
    SS14[39][22] = 4'h0;
    SS14[40][22] = 4'h0;
    SS14[41][22] = 4'h0;
    SS14[42][22] = 4'h0;
    SS14[43][22] = 4'h0;
    SS14[44][22] = 4'h0;
    SS14[45][22] = 4'h0;
    SS14[46][22] = 4'h0;
    SS14[47][22] = 4'h0;
    SS14[0][23] = 4'h0;
    SS14[1][23] = 4'h0;
    SS14[2][23] = 4'h0;
    SS14[3][23] = 4'h0;
    SS14[4][23] = 4'h0;
    SS14[5][23] = 4'h0;
    SS14[6][23] = 4'h0;
    SS14[7][23] = 4'h0;
    SS14[8][23] = 4'h0;
    SS14[9][23] = 4'h0;
    SS14[10][23] = 4'h0;
    SS14[11][23] = 4'h0;
    SS14[12][23] = 4'hD;
    SS14[13][23] = 4'hD;
    SS14[14][23] = 4'hD;
    SS14[15][23] = 4'hD;
    SS14[16][23] = 4'hD;
    SS14[17][23] = 4'hD;
    SS14[18][23] = 4'hC;
    SS14[19][23] = 4'hC;
    SS14[20][23] = 4'hC;
    SS14[21][23] = 4'hD;
    SS14[22][23] = 4'hD;
    SS14[23][23] = 4'hD;
    SS14[24][23] = 4'hD;
    SS14[25][23] = 4'hD;
    SS14[26][23] = 4'hD;
    SS14[27][23] = 4'hC;
    SS14[28][23] = 4'hC;
    SS14[29][23] = 4'hC;
    SS14[30][23] = 4'hD;
    SS14[31][23] = 4'hD;
    SS14[32][23] = 4'hD;
    SS14[33][23] = 4'hD;
    SS14[34][23] = 4'hD;
    SS14[35][23] = 4'hD;
    SS14[36][23] = 4'h0;
    SS14[37][23] = 4'h0;
    SS14[38][23] = 4'h0;
    SS14[39][23] = 4'h0;
    SS14[40][23] = 4'h0;
    SS14[41][23] = 4'h0;
    SS14[42][23] = 4'h0;
    SS14[43][23] = 4'h0;
    SS14[44][23] = 4'h0;
    SS14[45][23] = 4'h0;
    SS14[46][23] = 4'h0;
    SS14[47][23] = 4'h0;
    SS14[0][24] = 4'h0;
    SS14[1][24] = 4'h0;
    SS14[2][24] = 4'h0;
    SS14[3][24] = 4'h0;
    SS14[4][24] = 4'h0;
    SS14[5][24] = 4'h0;
    SS14[6][24] = 4'h3;
    SS14[7][24] = 4'h3;
    SS14[8][24] = 4'h3;
    SS14[9][24] = 4'hD;
    SS14[10][24] = 4'hD;
    SS14[11][24] = 4'hD;
    SS14[12][24] = 4'hD;
    SS14[13][24] = 4'hD;
    SS14[14][24] = 4'hD;
    SS14[15][24] = 4'hE;
    SS14[16][24] = 4'hE;
    SS14[17][24] = 4'hE;
    SS14[18][24] = 4'hC;
    SS14[19][24] = 4'hC;
    SS14[20][24] = 4'hC;
    SS14[21][24] = 4'hC;
    SS14[22][24] = 4'hC;
    SS14[23][24] = 4'hC;
    SS14[24][24] = 4'hC;
    SS14[25][24] = 4'hC;
    SS14[26][24] = 4'hC;
    SS14[27][24] = 4'hC;
    SS14[28][24] = 4'hC;
    SS14[29][24] = 4'hC;
    SS14[30][24] = 4'hE;
    SS14[31][24] = 4'hE;
    SS14[32][24] = 4'hE;
    SS14[33][24] = 4'hD;
    SS14[34][24] = 4'hD;
    SS14[35][24] = 4'hD;
    SS14[36][24] = 4'hD;
    SS14[37][24] = 4'hD;
    SS14[38][24] = 4'hD;
    SS14[39][24] = 4'h3;
    SS14[40][24] = 4'h3;
    SS14[41][24] = 4'h3;
    SS14[42][24] = 4'h0;
    SS14[43][24] = 4'h0;
    SS14[44][24] = 4'h0;
    SS14[45][24] = 4'h0;
    SS14[46][24] = 4'h0;
    SS14[47][24] = 4'h0;
    SS14[0][25] = 4'h0;
    SS14[1][25] = 4'h0;
    SS14[2][25] = 4'h0;
    SS14[3][25] = 4'h0;
    SS14[4][25] = 4'h0;
    SS14[5][25] = 4'h0;
    SS14[6][25] = 4'h3;
    SS14[7][25] = 4'h3;
    SS14[8][25] = 4'h3;
    SS14[9][25] = 4'hD;
    SS14[10][25] = 4'hD;
    SS14[11][25] = 4'hD;
    SS14[12][25] = 4'hD;
    SS14[13][25] = 4'hD;
    SS14[14][25] = 4'hD;
    SS14[15][25] = 4'hE;
    SS14[16][25] = 4'hE;
    SS14[17][25] = 4'hE;
    SS14[18][25] = 4'hC;
    SS14[19][25] = 4'hC;
    SS14[20][25] = 4'hC;
    SS14[21][25] = 4'hC;
    SS14[22][25] = 4'hC;
    SS14[23][25] = 4'hC;
    SS14[24][25] = 4'hC;
    SS14[25][25] = 4'hC;
    SS14[26][25] = 4'hC;
    SS14[27][25] = 4'hC;
    SS14[28][25] = 4'hC;
    SS14[29][25] = 4'hC;
    SS14[30][25] = 4'hE;
    SS14[31][25] = 4'hE;
    SS14[32][25] = 4'hE;
    SS14[33][25] = 4'hD;
    SS14[34][25] = 4'hD;
    SS14[35][25] = 4'hD;
    SS14[36][25] = 4'hD;
    SS14[37][25] = 4'hD;
    SS14[38][25] = 4'hD;
    SS14[39][25] = 4'h3;
    SS14[40][25] = 4'h3;
    SS14[41][25] = 4'h3;
    SS14[42][25] = 4'h0;
    SS14[43][25] = 4'h0;
    SS14[44][25] = 4'h0;
    SS14[45][25] = 4'h0;
    SS14[46][25] = 4'h0;
    SS14[47][25] = 4'h0;
    SS14[0][26] = 4'h0;
    SS14[1][26] = 4'h0;
    SS14[2][26] = 4'h0;
    SS14[3][26] = 4'h0;
    SS14[4][26] = 4'h0;
    SS14[5][26] = 4'h0;
    SS14[6][26] = 4'h3;
    SS14[7][26] = 4'h3;
    SS14[8][26] = 4'h3;
    SS14[9][26] = 4'hD;
    SS14[10][26] = 4'hD;
    SS14[11][26] = 4'hD;
    SS14[12][26] = 4'hD;
    SS14[13][26] = 4'hD;
    SS14[14][26] = 4'hD;
    SS14[15][26] = 4'hE;
    SS14[16][26] = 4'hE;
    SS14[17][26] = 4'hE;
    SS14[18][26] = 4'hC;
    SS14[19][26] = 4'hC;
    SS14[20][26] = 4'hC;
    SS14[21][26] = 4'hC;
    SS14[22][26] = 4'hC;
    SS14[23][26] = 4'hC;
    SS14[24][26] = 4'hC;
    SS14[25][26] = 4'hC;
    SS14[26][26] = 4'hC;
    SS14[27][26] = 4'hC;
    SS14[28][26] = 4'hC;
    SS14[29][26] = 4'hC;
    SS14[30][26] = 4'hE;
    SS14[31][26] = 4'hE;
    SS14[32][26] = 4'hE;
    SS14[33][26] = 4'hD;
    SS14[34][26] = 4'hD;
    SS14[35][26] = 4'hD;
    SS14[36][26] = 4'hD;
    SS14[37][26] = 4'hD;
    SS14[38][26] = 4'hD;
    SS14[39][26] = 4'h3;
    SS14[40][26] = 4'h3;
    SS14[41][26] = 4'h3;
    SS14[42][26] = 4'h0;
    SS14[43][26] = 4'h0;
    SS14[44][26] = 4'h0;
    SS14[45][26] = 4'h0;
    SS14[46][26] = 4'h0;
    SS14[47][26] = 4'h0;
    SS14[0][27] = 4'h0;
    SS14[1][27] = 4'h0;
    SS14[2][27] = 4'h0;
    SS14[3][27] = 4'hD;
    SS14[4][27] = 4'hD;
    SS14[5][27] = 4'hD;
    SS14[6][27] = 4'hD;
    SS14[7][27] = 4'hD;
    SS14[8][27] = 4'hD;
    SS14[9][27] = 4'hE;
    SS14[10][27] = 4'hE;
    SS14[11][27] = 4'hE;
    SS14[12][27] = 4'hE;
    SS14[13][27] = 4'hE;
    SS14[14][27] = 4'hE;
    SS14[15][27] = 4'hC;
    SS14[16][27] = 4'hC;
    SS14[17][27] = 4'hC;
    SS14[18][27] = 4'hC;
    SS14[19][27] = 4'hC;
    SS14[20][27] = 4'hC;
    SS14[21][27] = 4'hD;
    SS14[22][27] = 4'hD;
    SS14[23][27] = 4'hD;
    SS14[24][27] = 4'hD;
    SS14[25][27] = 4'hD;
    SS14[26][27] = 4'hD;
    SS14[27][27] = 4'hC;
    SS14[28][27] = 4'hC;
    SS14[29][27] = 4'hC;
    SS14[30][27] = 4'hC;
    SS14[31][27] = 4'hC;
    SS14[32][27] = 4'hC;
    SS14[33][27] = 4'hE;
    SS14[34][27] = 4'hE;
    SS14[35][27] = 4'hE;
    SS14[36][27] = 4'hE;
    SS14[37][27] = 4'hE;
    SS14[38][27] = 4'hE;
    SS14[39][27] = 4'hD;
    SS14[40][27] = 4'hD;
    SS14[41][27] = 4'hD;
    SS14[42][27] = 4'hD;
    SS14[43][27] = 4'hD;
    SS14[44][27] = 4'hD;
    SS14[45][27] = 4'h0;
    SS14[46][27] = 4'h0;
    SS14[47][27] = 4'h0;
    SS14[0][28] = 4'h0;
    SS14[1][28] = 4'h0;
    SS14[2][28] = 4'h0;
    SS14[3][28] = 4'hD;
    SS14[4][28] = 4'hD;
    SS14[5][28] = 4'hD;
    SS14[6][28] = 4'hD;
    SS14[7][28] = 4'hD;
    SS14[8][28] = 4'hD;
    SS14[9][28] = 4'hE;
    SS14[10][28] = 4'hE;
    SS14[11][28] = 4'hE;
    SS14[12][28] = 4'hE;
    SS14[13][28] = 4'hE;
    SS14[14][28] = 4'hE;
    SS14[15][28] = 4'hC;
    SS14[16][28] = 4'hC;
    SS14[17][28] = 4'hC;
    SS14[18][28] = 4'hC;
    SS14[19][28] = 4'hC;
    SS14[20][28] = 4'hC;
    SS14[21][28] = 4'hD;
    SS14[22][28] = 4'hD;
    SS14[23][28] = 4'hD;
    SS14[24][28] = 4'hD;
    SS14[25][28] = 4'hD;
    SS14[26][28] = 4'hD;
    SS14[27][28] = 4'hC;
    SS14[28][28] = 4'hC;
    SS14[29][28] = 4'hC;
    SS14[30][28] = 4'hC;
    SS14[31][28] = 4'hC;
    SS14[32][28] = 4'hC;
    SS14[33][28] = 4'hE;
    SS14[34][28] = 4'hE;
    SS14[35][28] = 4'hE;
    SS14[36][28] = 4'hE;
    SS14[37][28] = 4'hE;
    SS14[38][28] = 4'hE;
    SS14[39][28] = 4'hD;
    SS14[40][28] = 4'hD;
    SS14[41][28] = 4'hD;
    SS14[42][28] = 4'hD;
    SS14[43][28] = 4'hD;
    SS14[44][28] = 4'hD;
    SS14[45][28] = 4'h0;
    SS14[46][28] = 4'h0;
    SS14[47][28] = 4'h0;
    SS14[0][29] = 4'h0;
    SS14[1][29] = 4'h0;
    SS14[2][29] = 4'h0;
    SS14[3][29] = 4'hD;
    SS14[4][29] = 4'hD;
    SS14[5][29] = 4'hD;
    SS14[6][29] = 4'hD;
    SS14[7][29] = 4'hD;
    SS14[8][29] = 4'hD;
    SS14[9][29] = 4'hE;
    SS14[10][29] = 4'hE;
    SS14[11][29] = 4'hE;
    SS14[12][29] = 4'hE;
    SS14[13][29] = 4'hE;
    SS14[14][29] = 4'hE;
    SS14[15][29] = 4'hC;
    SS14[16][29] = 4'hC;
    SS14[17][29] = 4'hC;
    SS14[18][29] = 4'hC;
    SS14[19][29] = 4'hC;
    SS14[20][29] = 4'hC;
    SS14[21][29] = 4'hD;
    SS14[22][29] = 4'hD;
    SS14[23][29] = 4'hD;
    SS14[24][29] = 4'hD;
    SS14[25][29] = 4'hD;
    SS14[26][29] = 4'hD;
    SS14[27][29] = 4'hC;
    SS14[28][29] = 4'hC;
    SS14[29][29] = 4'hC;
    SS14[30][29] = 4'hC;
    SS14[31][29] = 4'hC;
    SS14[32][29] = 4'hC;
    SS14[33][29] = 4'hE;
    SS14[34][29] = 4'hE;
    SS14[35][29] = 4'hE;
    SS14[36][29] = 4'hE;
    SS14[37][29] = 4'hE;
    SS14[38][29] = 4'hE;
    SS14[39][29] = 4'hD;
    SS14[40][29] = 4'hD;
    SS14[41][29] = 4'hD;
    SS14[42][29] = 4'hD;
    SS14[43][29] = 4'hD;
    SS14[44][29] = 4'hD;
    SS14[45][29] = 4'h0;
    SS14[46][29] = 4'h0;
    SS14[47][29] = 4'h0;
    SS14[0][30] = 4'hD;
    SS14[1][30] = 4'hD;
    SS14[2][30] = 4'hD;
    SS14[3][30] = 4'hD;
    SS14[4][30] = 4'hD;
    SS14[5][30] = 4'hD;
    SS14[6][30] = 4'hE;
    SS14[7][30] = 4'hE;
    SS14[8][30] = 4'hE;
    SS14[9][30] = 4'hE;
    SS14[10][30] = 4'hE;
    SS14[11][30] = 4'hE;
    SS14[12][30] = 4'hC;
    SS14[13][30] = 4'hC;
    SS14[14][30] = 4'hC;
    SS14[15][30] = 4'hC;
    SS14[16][30] = 4'hC;
    SS14[17][30] = 4'hC;
    SS14[18][30] = 4'hC;
    SS14[19][30] = 4'hC;
    SS14[20][30] = 4'hC;
    SS14[21][30] = 4'hE;
    SS14[22][30] = 4'hE;
    SS14[23][30] = 4'hE;
    SS14[24][30] = 4'hE;
    SS14[25][30] = 4'hE;
    SS14[26][30] = 4'hE;
    SS14[27][30] = 4'hC;
    SS14[28][30] = 4'hC;
    SS14[29][30] = 4'hC;
    SS14[30][30] = 4'hC;
    SS14[31][30] = 4'hC;
    SS14[32][30] = 4'hC;
    SS14[33][30] = 4'hC;
    SS14[34][30] = 4'hC;
    SS14[35][30] = 4'hC;
    SS14[36][30] = 4'hE;
    SS14[37][30] = 4'hE;
    SS14[38][30] = 4'hE;
    SS14[39][30] = 4'hE;
    SS14[40][30] = 4'hE;
    SS14[41][30] = 4'hE;
    SS14[42][30] = 4'hD;
    SS14[43][30] = 4'hD;
    SS14[44][30] = 4'hD;
    SS14[45][30] = 4'hD;
    SS14[46][30] = 4'hD;
    SS14[47][30] = 4'hD;
    SS14[0][31] = 4'hD;
    SS14[1][31] = 4'hD;
    SS14[2][31] = 4'hD;
    SS14[3][31] = 4'hD;
    SS14[4][31] = 4'hD;
    SS14[5][31] = 4'hD;
    SS14[6][31] = 4'hE;
    SS14[7][31] = 4'hE;
    SS14[8][31] = 4'hE;
    SS14[9][31] = 4'hE;
    SS14[10][31] = 4'hE;
    SS14[11][31] = 4'hE;
    SS14[12][31] = 4'hC;
    SS14[13][31] = 4'hC;
    SS14[14][31] = 4'hC;
    SS14[15][31] = 4'hC;
    SS14[16][31] = 4'hC;
    SS14[17][31] = 4'hC;
    SS14[18][31] = 4'hC;
    SS14[19][31] = 4'hC;
    SS14[20][31] = 4'hC;
    SS14[21][31] = 4'hE;
    SS14[22][31] = 4'hE;
    SS14[23][31] = 4'hE;
    SS14[24][31] = 4'hE;
    SS14[25][31] = 4'hE;
    SS14[26][31] = 4'hE;
    SS14[27][31] = 4'hC;
    SS14[28][31] = 4'hC;
    SS14[29][31] = 4'hC;
    SS14[30][31] = 4'hC;
    SS14[31][31] = 4'hC;
    SS14[32][31] = 4'hC;
    SS14[33][31] = 4'hC;
    SS14[34][31] = 4'hC;
    SS14[35][31] = 4'hC;
    SS14[36][31] = 4'hE;
    SS14[37][31] = 4'hE;
    SS14[38][31] = 4'hE;
    SS14[39][31] = 4'hE;
    SS14[40][31] = 4'hE;
    SS14[41][31] = 4'hE;
    SS14[42][31] = 4'hD;
    SS14[43][31] = 4'hD;
    SS14[44][31] = 4'hD;
    SS14[45][31] = 4'hD;
    SS14[46][31] = 4'hD;
    SS14[47][31] = 4'hD;
    SS14[0][32] = 4'hD;
    SS14[1][32] = 4'hD;
    SS14[2][32] = 4'hD;
    SS14[3][32] = 4'hD;
    SS14[4][32] = 4'hD;
    SS14[5][32] = 4'hD;
    SS14[6][32] = 4'hE;
    SS14[7][32] = 4'hE;
    SS14[8][32] = 4'hE;
    SS14[9][32] = 4'hE;
    SS14[10][32] = 4'hE;
    SS14[11][32] = 4'hE;
    SS14[12][32] = 4'hC;
    SS14[13][32] = 4'hC;
    SS14[14][32] = 4'hC;
    SS14[15][32] = 4'hC;
    SS14[16][32] = 4'hC;
    SS14[17][32] = 4'hC;
    SS14[18][32] = 4'hC;
    SS14[19][32] = 4'hC;
    SS14[20][32] = 4'hC;
    SS14[21][32] = 4'hE;
    SS14[22][32] = 4'hE;
    SS14[23][32] = 4'hE;
    SS14[24][32] = 4'hE;
    SS14[25][32] = 4'hE;
    SS14[26][32] = 4'hE;
    SS14[27][32] = 4'hC;
    SS14[28][32] = 4'hC;
    SS14[29][32] = 4'hC;
    SS14[30][32] = 4'hC;
    SS14[31][32] = 4'hC;
    SS14[32][32] = 4'hC;
    SS14[33][32] = 4'hC;
    SS14[34][32] = 4'hC;
    SS14[35][32] = 4'hC;
    SS14[36][32] = 4'hE;
    SS14[37][32] = 4'hE;
    SS14[38][32] = 4'hE;
    SS14[39][32] = 4'hE;
    SS14[40][32] = 4'hE;
    SS14[41][32] = 4'hE;
    SS14[42][32] = 4'hD;
    SS14[43][32] = 4'hD;
    SS14[44][32] = 4'hD;
    SS14[45][32] = 4'hD;
    SS14[46][32] = 4'hD;
    SS14[47][32] = 4'hD;
    SS14[0][33] = 4'h0;
    SS14[1][33] = 4'h0;
    SS14[2][33] = 4'h0;
    SS14[3][33] = 4'h0;
    SS14[4][33] = 4'h0;
    SS14[5][33] = 4'h0;
    SS14[6][33] = 4'h0;
    SS14[7][33] = 4'h0;
    SS14[8][33] = 4'h0;
    SS14[9][33] = 4'h0;
    SS14[10][33] = 4'h0;
    SS14[11][33] = 4'h0;
    SS14[12][33] = 4'hC;
    SS14[13][33] = 4'hC;
    SS14[14][33] = 4'hC;
    SS14[15][33] = 4'hC;
    SS14[16][33] = 4'hC;
    SS14[17][33] = 4'hC;
    SS14[18][33] = 4'hD;
    SS14[19][33] = 4'hD;
    SS14[20][33] = 4'hD;
    SS14[21][33] = 4'hE;
    SS14[22][33] = 4'hE;
    SS14[23][33] = 4'hE;
    SS14[24][33] = 4'hE;
    SS14[25][33] = 4'hE;
    SS14[26][33] = 4'hE;
    SS14[27][33] = 4'hD;
    SS14[28][33] = 4'hD;
    SS14[29][33] = 4'hD;
    SS14[30][33] = 4'hC;
    SS14[31][33] = 4'hC;
    SS14[32][33] = 4'hC;
    SS14[33][33] = 4'hC;
    SS14[34][33] = 4'hC;
    SS14[35][33] = 4'hC;
    SS14[36][33] = 4'h0;
    SS14[37][33] = 4'h0;
    SS14[38][33] = 4'h0;
    SS14[39][33] = 4'h0;
    SS14[40][33] = 4'h0;
    SS14[41][33] = 4'h0;
    SS14[42][33] = 4'h0;
    SS14[43][33] = 4'h0;
    SS14[44][33] = 4'h0;
    SS14[45][33] = 4'h0;
    SS14[46][33] = 4'h0;
    SS14[47][33] = 4'h0;
    SS14[0][34] = 4'h0;
    SS14[1][34] = 4'h0;
    SS14[2][34] = 4'h0;
    SS14[3][34] = 4'h0;
    SS14[4][34] = 4'h0;
    SS14[5][34] = 4'h0;
    SS14[6][34] = 4'h0;
    SS14[7][34] = 4'h0;
    SS14[8][34] = 4'h0;
    SS14[9][34] = 4'h0;
    SS14[10][34] = 4'h0;
    SS14[11][34] = 4'h0;
    SS14[12][34] = 4'hC;
    SS14[13][34] = 4'hC;
    SS14[14][34] = 4'hC;
    SS14[15][34] = 4'hC;
    SS14[16][34] = 4'hC;
    SS14[17][34] = 4'hC;
    SS14[18][34] = 4'hD;
    SS14[19][34] = 4'hD;
    SS14[20][34] = 4'hD;
    SS14[21][34] = 4'hE;
    SS14[22][34] = 4'hE;
    SS14[23][34] = 4'hE;
    SS14[24][34] = 4'hE;
    SS14[25][34] = 4'hE;
    SS14[26][34] = 4'hE;
    SS14[27][34] = 4'hD;
    SS14[28][34] = 4'hD;
    SS14[29][34] = 4'hD;
    SS14[30][34] = 4'hC;
    SS14[31][34] = 4'hC;
    SS14[32][34] = 4'hC;
    SS14[33][34] = 4'hC;
    SS14[34][34] = 4'hC;
    SS14[35][34] = 4'hC;
    SS14[36][34] = 4'h0;
    SS14[37][34] = 4'h0;
    SS14[38][34] = 4'h0;
    SS14[39][34] = 4'h0;
    SS14[40][34] = 4'h0;
    SS14[41][34] = 4'h0;
    SS14[42][34] = 4'h0;
    SS14[43][34] = 4'h0;
    SS14[44][34] = 4'h0;
    SS14[45][34] = 4'h0;
    SS14[46][34] = 4'h0;
    SS14[47][34] = 4'h0;
    SS14[0][35] = 4'h0;
    SS14[1][35] = 4'h0;
    SS14[2][35] = 4'h0;
    SS14[3][35] = 4'h0;
    SS14[4][35] = 4'h0;
    SS14[5][35] = 4'h0;
    SS14[6][35] = 4'h0;
    SS14[7][35] = 4'h0;
    SS14[8][35] = 4'h0;
    SS14[9][35] = 4'h0;
    SS14[10][35] = 4'h0;
    SS14[11][35] = 4'h0;
    SS14[12][35] = 4'hC;
    SS14[13][35] = 4'hC;
    SS14[14][35] = 4'hC;
    SS14[15][35] = 4'hC;
    SS14[16][35] = 4'hC;
    SS14[17][35] = 4'hC;
    SS14[18][35] = 4'hD;
    SS14[19][35] = 4'hD;
    SS14[20][35] = 4'hD;
    SS14[21][35] = 4'hE;
    SS14[22][35] = 4'hE;
    SS14[23][35] = 4'hE;
    SS14[24][35] = 4'hE;
    SS14[25][35] = 4'hE;
    SS14[26][35] = 4'hE;
    SS14[27][35] = 4'hD;
    SS14[28][35] = 4'hD;
    SS14[29][35] = 4'hD;
    SS14[30][35] = 4'hC;
    SS14[31][35] = 4'hC;
    SS14[32][35] = 4'hC;
    SS14[33][35] = 4'hC;
    SS14[34][35] = 4'hC;
    SS14[35][35] = 4'hC;
    SS14[36][35] = 4'h0;
    SS14[37][35] = 4'h0;
    SS14[38][35] = 4'h0;
    SS14[39][35] = 4'h0;
    SS14[40][35] = 4'h0;
    SS14[41][35] = 4'h0;
    SS14[42][35] = 4'h0;
    SS14[43][35] = 4'h0;
    SS14[44][35] = 4'h0;
    SS14[45][35] = 4'h0;
    SS14[46][35] = 4'h0;
    SS14[47][35] = 4'h0;
    SS14[0][36] = 4'h0;
    SS14[1][36] = 4'h0;
    SS14[2][36] = 4'h0;
    SS14[3][36] = 4'h0;
    SS14[4][36] = 4'h0;
    SS14[5][36] = 4'h0;
    SS14[6][36] = 4'h0;
    SS14[7][36] = 4'h0;
    SS14[8][36] = 4'h0;
    SS14[9][36] = 4'h0;
    SS14[10][36] = 4'h0;
    SS14[11][36] = 4'h0;
    SS14[12][36] = 4'hC;
    SS14[13][36] = 4'hC;
    SS14[14][36] = 4'hC;
    SS14[15][36] = 4'hD;
    SS14[16][36] = 4'hD;
    SS14[17][36] = 4'hD;
    SS14[18][36] = 4'hE;
    SS14[19][36] = 4'hE;
    SS14[20][36] = 4'hE;
    SS14[21][36] = 4'h0;
    SS14[22][36] = 4'h0;
    SS14[23][36] = 4'h0;
    SS14[24][36] = 4'h0;
    SS14[25][36] = 4'h0;
    SS14[26][36] = 4'h0;
    SS14[27][36] = 4'hE;
    SS14[28][36] = 4'hE;
    SS14[29][36] = 4'hE;
    SS14[30][36] = 4'hD;
    SS14[31][36] = 4'hD;
    SS14[32][36] = 4'hD;
    SS14[33][36] = 4'hC;
    SS14[34][36] = 4'hC;
    SS14[35][36] = 4'hC;
    SS14[36][36] = 4'h0;
    SS14[37][36] = 4'h0;
    SS14[38][36] = 4'h0;
    SS14[39][36] = 4'h0;
    SS14[40][36] = 4'h0;
    SS14[41][36] = 4'h0;
    SS14[42][36] = 4'h0;
    SS14[43][36] = 4'h0;
    SS14[44][36] = 4'h0;
    SS14[45][36] = 4'h0;
    SS14[46][36] = 4'h0;
    SS14[47][36] = 4'h0;
    SS14[0][37] = 4'h0;
    SS14[1][37] = 4'h0;
    SS14[2][37] = 4'h0;
    SS14[3][37] = 4'h0;
    SS14[4][37] = 4'h0;
    SS14[5][37] = 4'h0;
    SS14[6][37] = 4'h0;
    SS14[7][37] = 4'h0;
    SS14[8][37] = 4'h0;
    SS14[9][37] = 4'h0;
    SS14[10][37] = 4'h0;
    SS14[11][37] = 4'h0;
    SS14[12][37] = 4'hC;
    SS14[13][37] = 4'hC;
    SS14[14][37] = 4'hC;
    SS14[15][37] = 4'hD;
    SS14[16][37] = 4'hD;
    SS14[17][37] = 4'hD;
    SS14[18][37] = 4'hE;
    SS14[19][37] = 4'hE;
    SS14[20][37] = 4'hE;
    SS14[21][37] = 4'h0;
    SS14[22][37] = 4'h0;
    SS14[23][37] = 4'h0;
    SS14[24][37] = 4'h0;
    SS14[25][37] = 4'h0;
    SS14[26][37] = 4'h0;
    SS14[27][37] = 4'hE;
    SS14[28][37] = 4'hE;
    SS14[29][37] = 4'hE;
    SS14[30][37] = 4'hD;
    SS14[31][37] = 4'hD;
    SS14[32][37] = 4'hD;
    SS14[33][37] = 4'hC;
    SS14[34][37] = 4'hC;
    SS14[35][37] = 4'hC;
    SS14[36][37] = 4'h0;
    SS14[37][37] = 4'h0;
    SS14[38][37] = 4'h0;
    SS14[39][37] = 4'h0;
    SS14[40][37] = 4'h0;
    SS14[41][37] = 4'h0;
    SS14[42][37] = 4'h0;
    SS14[43][37] = 4'h0;
    SS14[44][37] = 4'h0;
    SS14[45][37] = 4'h0;
    SS14[46][37] = 4'h0;
    SS14[47][37] = 4'h0;
    SS14[0][38] = 4'h0;
    SS14[1][38] = 4'h0;
    SS14[2][38] = 4'h0;
    SS14[3][38] = 4'h0;
    SS14[4][38] = 4'h0;
    SS14[5][38] = 4'h0;
    SS14[6][38] = 4'h0;
    SS14[7][38] = 4'h0;
    SS14[8][38] = 4'h0;
    SS14[9][38] = 4'h0;
    SS14[10][38] = 4'h0;
    SS14[11][38] = 4'h0;
    SS14[12][38] = 4'hC;
    SS14[13][38] = 4'hC;
    SS14[14][38] = 4'hC;
    SS14[15][38] = 4'hD;
    SS14[16][38] = 4'hD;
    SS14[17][38] = 4'hD;
    SS14[18][38] = 4'hE;
    SS14[19][38] = 4'hE;
    SS14[20][38] = 4'hE;
    SS14[21][38] = 4'h0;
    SS14[22][38] = 4'h0;
    SS14[23][38] = 4'h0;
    SS14[24][38] = 4'h0;
    SS14[25][38] = 4'h0;
    SS14[26][38] = 4'h0;
    SS14[27][38] = 4'hE;
    SS14[28][38] = 4'hE;
    SS14[29][38] = 4'hE;
    SS14[30][38] = 4'hD;
    SS14[31][38] = 4'hD;
    SS14[32][38] = 4'hD;
    SS14[33][38] = 4'hC;
    SS14[34][38] = 4'hC;
    SS14[35][38] = 4'hC;
    SS14[36][38] = 4'h0;
    SS14[37][38] = 4'h0;
    SS14[38][38] = 4'h0;
    SS14[39][38] = 4'h0;
    SS14[40][38] = 4'h0;
    SS14[41][38] = 4'h0;
    SS14[42][38] = 4'h0;
    SS14[43][38] = 4'h0;
    SS14[44][38] = 4'h0;
    SS14[45][38] = 4'h0;
    SS14[46][38] = 4'h0;
    SS14[47][38] = 4'h0;
    SS14[0][39] = 4'h0;
    SS14[1][39] = 4'h0;
    SS14[2][39] = 4'h0;
    SS14[3][39] = 4'h0;
    SS14[4][39] = 4'h0;
    SS14[5][39] = 4'h0;
    SS14[6][39] = 4'h0;
    SS14[7][39] = 4'h0;
    SS14[8][39] = 4'h0;
    SS14[9][39] = 4'hC;
    SS14[10][39] = 4'hC;
    SS14[11][39] = 4'hC;
    SS14[12][39] = 4'hC;
    SS14[13][39] = 4'hC;
    SS14[14][39] = 4'hC;
    SS14[15][39] = 4'hE;
    SS14[16][39] = 4'hE;
    SS14[17][39] = 4'hE;
    SS14[18][39] = 4'h0;
    SS14[19][39] = 4'h0;
    SS14[20][39] = 4'h0;
    SS14[21][39] = 4'h0;
    SS14[22][39] = 4'h0;
    SS14[23][39] = 4'h0;
    SS14[24][39] = 4'h0;
    SS14[25][39] = 4'h0;
    SS14[26][39] = 4'h0;
    SS14[27][39] = 4'h0;
    SS14[28][39] = 4'h0;
    SS14[29][39] = 4'h0;
    SS14[30][39] = 4'hE;
    SS14[31][39] = 4'hE;
    SS14[32][39] = 4'hE;
    SS14[33][39] = 4'hC;
    SS14[34][39] = 4'hC;
    SS14[35][39] = 4'hC;
    SS14[36][39] = 4'hC;
    SS14[37][39] = 4'hC;
    SS14[38][39] = 4'hC;
    SS14[39][39] = 4'h0;
    SS14[40][39] = 4'h0;
    SS14[41][39] = 4'h0;
    SS14[42][39] = 4'h0;
    SS14[43][39] = 4'h0;
    SS14[44][39] = 4'h0;
    SS14[45][39] = 4'h0;
    SS14[46][39] = 4'h0;
    SS14[47][39] = 4'h0;
    SS14[0][40] = 4'h0;
    SS14[1][40] = 4'h0;
    SS14[2][40] = 4'h0;
    SS14[3][40] = 4'h0;
    SS14[4][40] = 4'h0;
    SS14[5][40] = 4'h0;
    SS14[6][40] = 4'h0;
    SS14[7][40] = 4'h0;
    SS14[8][40] = 4'h0;
    SS14[9][40] = 4'hC;
    SS14[10][40] = 4'hC;
    SS14[11][40] = 4'hC;
    SS14[12][40] = 4'hC;
    SS14[13][40] = 4'hC;
    SS14[14][40] = 4'hC;
    SS14[15][40] = 4'hE;
    SS14[16][40] = 4'hE;
    SS14[17][40] = 4'hE;
    SS14[18][40] = 4'h0;
    SS14[19][40] = 4'h0;
    SS14[20][40] = 4'h0;
    SS14[21][40] = 4'h0;
    SS14[22][40] = 4'h0;
    SS14[23][40] = 4'h0;
    SS14[24][40] = 4'h0;
    SS14[25][40] = 4'h0;
    SS14[26][40] = 4'h0;
    SS14[27][40] = 4'h0;
    SS14[28][40] = 4'h0;
    SS14[29][40] = 4'h0;
    SS14[30][40] = 4'hE;
    SS14[31][40] = 4'hE;
    SS14[32][40] = 4'hE;
    SS14[33][40] = 4'hC;
    SS14[34][40] = 4'hC;
    SS14[35][40] = 4'hC;
    SS14[36][40] = 4'hC;
    SS14[37][40] = 4'hC;
    SS14[38][40] = 4'hC;
    SS14[39][40] = 4'h0;
    SS14[40][40] = 4'h0;
    SS14[41][40] = 4'h0;
    SS14[42][40] = 4'h0;
    SS14[43][40] = 4'h0;
    SS14[44][40] = 4'h0;
    SS14[45][40] = 4'h0;
    SS14[46][40] = 4'h0;
    SS14[47][40] = 4'h0;
    SS14[0][41] = 4'h0;
    SS14[1][41] = 4'h0;
    SS14[2][41] = 4'h0;
    SS14[3][41] = 4'h0;
    SS14[4][41] = 4'h0;
    SS14[5][41] = 4'h0;
    SS14[6][41] = 4'h0;
    SS14[7][41] = 4'h0;
    SS14[8][41] = 4'h0;
    SS14[9][41] = 4'hC;
    SS14[10][41] = 4'hC;
    SS14[11][41] = 4'hC;
    SS14[12][41] = 4'hC;
    SS14[13][41] = 4'hC;
    SS14[14][41] = 4'hC;
    SS14[15][41] = 4'hE;
    SS14[16][41] = 4'hE;
    SS14[17][41] = 4'hE;
    SS14[18][41] = 4'h0;
    SS14[19][41] = 4'h0;
    SS14[20][41] = 4'h0;
    SS14[21][41] = 4'h0;
    SS14[22][41] = 4'h0;
    SS14[23][41] = 4'h0;
    SS14[24][41] = 4'h0;
    SS14[25][41] = 4'h0;
    SS14[26][41] = 4'h0;
    SS14[27][41] = 4'h0;
    SS14[28][41] = 4'h0;
    SS14[29][41] = 4'h0;
    SS14[30][41] = 4'hE;
    SS14[31][41] = 4'hE;
    SS14[32][41] = 4'hE;
    SS14[33][41] = 4'hC;
    SS14[34][41] = 4'hC;
    SS14[35][41] = 4'hC;
    SS14[36][41] = 4'hC;
    SS14[37][41] = 4'hC;
    SS14[38][41] = 4'hC;
    SS14[39][41] = 4'h0;
    SS14[40][41] = 4'h0;
    SS14[41][41] = 4'h0;
    SS14[42][41] = 4'h0;
    SS14[43][41] = 4'h0;
    SS14[44][41] = 4'h0;
    SS14[45][41] = 4'h0;
    SS14[46][41] = 4'h0;
    SS14[47][41] = 4'h0;
    SS14[0][42] = 4'h0;
    SS14[1][42] = 4'h0;
    SS14[2][42] = 4'h0;
    SS14[3][42] = 4'h0;
    SS14[4][42] = 4'h0;
    SS14[5][42] = 4'h0;
    SS14[6][42] = 4'h0;
    SS14[7][42] = 4'h0;
    SS14[8][42] = 4'h0;
    SS14[9][42] = 4'hC;
    SS14[10][42] = 4'hC;
    SS14[11][42] = 4'hC;
    SS14[12][42] = 4'hD;
    SS14[13][42] = 4'hD;
    SS14[14][42] = 4'hD;
    SS14[15][42] = 4'h0;
    SS14[16][42] = 4'h0;
    SS14[17][42] = 4'h0;
    SS14[18][42] = 4'h0;
    SS14[19][42] = 4'h0;
    SS14[20][42] = 4'h0;
    SS14[21][42] = 4'h0;
    SS14[22][42] = 4'h0;
    SS14[23][42] = 4'h0;
    SS14[24][42] = 4'h0;
    SS14[25][42] = 4'h0;
    SS14[26][42] = 4'h0;
    SS14[27][42] = 4'h0;
    SS14[28][42] = 4'h0;
    SS14[29][42] = 4'h0;
    SS14[30][42] = 4'h0;
    SS14[31][42] = 4'h0;
    SS14[32][42] = 4'h0;
    SS14[33][42] = 4'hD;
    SS14[34][42] = 4'hD;
    SS14[35][42] = 4'hD;
    SS14[36][42] = 4'hC;
    SS14[37][42] = 4'hC;
    SS14[38][42] = 4'hC;
    SS14[39][42] = 4'h0;
    SS14[40][42] = 4'h0;
    SS14[41][42] = 4'h0;
    SS14[42][42] = 4'h0;
    SS14[43][42] = 4'h0;
    SS14[44][42] = 4'h0;
    SS14[45][42] = 4'h0;
    SS14[46][42] = 4'h0;
    SS14[47][42] = 4'h0;
    SS14[0][43] = 4'h0;
    SS14[1][43] = 4'h0;
    SS14[2][43] = 4'h0;
    SS14[3][43] = 4'h0;
    SS14[4][43] = 4'h0;
    SS14[5][43] = 4'h0;
    SS14[6][43] = 4'h0;
    SS14[7][43] = 4'h0;
    SS14[8][43] = 4'h0;
    SS14[9][43] = 4'hC;
    SS14[10][43] = 4'hC;
    SS14[11][43] = 4'hC;
    SS14[12][43] = 4'hD;
    SS14[13][43] = 4'hD;
    SS14[14][43] = 4'hD;
    SS14[15][43] = 4'h0;
    SS14[16][43] = 4'h0;
    SS14[17][43] = 4'h0;
    SS14[18][43] = 4'h0;
    SS14[19][43] = 4'h0;
    SS14[20][43] = 4'h0;
    SS14[21][43] = 4'h0;
    SS14[22][43] = 4'h0;
    SS14[23][43] = 4'h0;
    SS14[24][43] = 4'h0;
    SS14[25][43] = 4'h0;
    SS14[26][43] = 4'h0;
    SS14[27][43] = 4'h0;
    SS14[28][43] = 4'h0;
    SS14[29][43] = 4'h0;
    SS14[30][43] = 4'h0;
    SS14[31][43] = 4'h0;
    SS14[32][43] = 4'h0;
    SS14[33][43] = 4'hD;
    SS14[34][43] = 4'hD;
    SS14[35][43] = 4'hD;
    SS14[36][43] = 4'hC;
    SS14[37][43] = 4'hC;
    SS14[38][43] = 4'hC;
    SS14[39][43] = 4'h0;
    SS14[40][43] = 4'h0;
    SS14[41][43] = 4'h0;
    SS14[42][43] = 4'h0;
    SS14[43][43] = 4'h0;
    SS14[44][43] = 4'h0;
    SS14[45][43] = 4'h0;
    SS14[46][43] = 4'h0;
    SS14[47][43] = 4'h0;
    SS14[0][44] = 4'h0;
    SS14[1][44] = 4'h0;
    SS14[2][44] = 4'h0;
    SS14[3][44] = 4'h0;
    SS14[4][44] = 4'h0;
    SS14[5][44] = 4'h0;
    SS14[6][44] = 4'h0;
    SS14[7][44] = 4'h0;
    SS14[8][44] = 4'h0;
    SS14[9][44] = 4'hC;
    SS14[10][44] = 4'hC;
    SS14[11][44] = 4'hC;
    SS14[12][44] = 4'hD;
    SS14[13][44] = 4'hD;
    SS14[14][44] = 4'hD;
    SS14[15][44] = 4'h0;
    SS14[16][44] = 4'h0;
    SS14[17][44] = 4'h0;
    SS14[18][44] = 4'h0;
    SS14[19][44] = 4'h0;
    SS14[20][44] = 4'h0;
    SS14[21][44] = 4'h0;
    SS14[22][44] = 4'h0;
    SS14[23][44] = 4'h0;
    SS14[24][44] = 4'h0;
    SS14[25][44] = 4'h0;
    SS14[26][44] = 4'h0;
    SS14[27][44] = 4'h0;
    SS14[28][44] = 4'h0;
    SS14[29][44] = 4'h0;
    SS14[30][44] = 4'h0;
    SS14[31][44] = 4'h0;
    SS14[32][44] = 4'h0;
    SS14[33][44] = 4'hD;
    SS14[34][44] = 4'hD;
    SS14[35][44] = 4'hD;
    SS14[36][44] = 4'hC;
    SS14[37][44] = 4'hC;
    SS14[38][44] = 4'hC;
    SS14[39][44] = 4'h0;
    SS14[40][44] = 4'h0;
    SS14[41][44] = 4'h0;
    SS14[42][44] = 4'h0;
    SS14[43][44] = 4'h0;
    SS14[44][44] = 4'h0;
    SS14[45][44] = 4'h0;
    SS14[46][44] = 4'h0;
    SS14[47][44] = 4'h0;
    SS14[0][45] = 4'h0;
    SS14[1][45] = 4'h0;
    SS14[2][45] = 4'h0;
    SS14[3][45] = 4'h0;
    SS14[4][45] = 4'h0;
    SS14[5][45] = 4'h0;
    SS14[6][45] = 4'h0;
    SS14[7][45] = 4'h0;
    SS14[8][45] = 4'h0;
    SS14[9][45] = 4'hD;
    SS14[10][45] = 4'hD;
    SS14[11][45] = 4'hD;
    SS14[12][45] = 4'h0;
    SS14[13][45] = 4'h0;
    SS14[14][45] = 4'h0;
    SS14[15][45] = 4'h0;
    SS14[16][45] = 4'h0;
    SS14[17][45] = 4'h0;
    SS14[18][45] = 4'h0;
    SS14[19][45] = 4'h0;
    SS14[20][45] = 4'h0;
    SS14[21][45] = 4'h0;
    SS14[22][45] = 4'h0;
    SS14[23][45] = 4'h0;
    SS14[24][45] = 4'h0;
    SS14[25][45] = 4'h0;
    SS14[26][45] = 4'h0;
    SS14[27][45] = 4'h0;
    SS14[28][45] = 4'h0;
    SS14[29][45] = 4'h0;
    SS14[30][45] = 4'h0;
    SS14[31][45] = 4'h0;
    SS14[32][45] = 4'h0;
    SS14[33][45] = 4'h0;
    SS14[34][45] = 4'h0;
    SS14[35][45] = 4'h0;
    SS14[36][45] = 4'hD;
    SS14[37][45] = 4'hD;
    SS14[38][45] = 4'hD;
    SS14[39][45] = 4'h0;
    SS14[40][45] = 4'h0;
    SS14[41][45] = 4'h0;
    SS14[42][45] = 4'h0;
    SS14[43][45] = 4'h0;
    SS14[44][45] = 4'h0;
    SS14[45][45] = 4'h0;
    SS14[46][45] = 4'h0;
    SS14[47][45] = 4'h0;
    SS14[0][46] = 4'h0;
    SS14[1][46] = 4'h0;
    SS14[2][46] = 4'h0;
    SS14[3][46] = 4'h0;
    SS14[4][46] = 4'h0;
    SS14[5][46] = 4'h0;
    SS14[6][46] = 4'h0;
    SS14[7][46] = 4'h0;
    SS14[8][46] = 4'h0;
    SS14[9][46] = 4'hD;
    SS14[10][46] = 4'hD;
    SS14[11][46] = 4'hD;
    SS14[12][46] = 4'h0;
    SS14[13][46] = 4'h0;
    SS14[14][46] = 4'h0;
    SS14[15][46] = 4'h0;
    SS14[16][46] = 4'h0;
    SS14[17][46] = 4'h0;
    SS14[18][46] = 4'h0;
    SS14[19][46] = 4'h0;
    SS14[20][46] = 4'h0;
    SS14[21][46] = 4'h0;
    SS14[22][46] = 4'h0;
    SS14[23][46] = 4'h0;
    SS14[24][46] = 4'h0;
    SS14[25][46] = 4'h0;
    SS14[26][46] = 4'h0;
    SS14[27][46] = 4'h0;
    SS14[28][46] = 4'h0;
    SS14[29][46] = 4'h0;
    SS14[30][46] = 4'h0;
    SS14[31][46] = 4'h0;
    SS14[32][46] = 4'h0;
    SS14[33][46] = 4'h0;
    SS14[34][46] = 4'h0;
    SS14[35][46] = 4'h0;
    SS14[36][46] = 4'hD;
    SS14[37][46] = 4'hD;
    SS14[38][46] = 4'hD;
    SS14[39][46] = 4'h0;
    SS14[40][46] = 4'h0;
    SS14[41][46] = 4'h0;
    SS14[42][46] = 4'h0;
    SS14[43][46] = 4'h0;
    SS14[44][46] = 4'h0;
    SS14[45][46] = 4'h0;
    SS14[46][46] = 4'h0;
    SS14[47][46] = 4'h0;
    SS14[0][47] = 4'h0;
    SS14[1][47] = 4'h0;
    SS14[2][47] = 4'h0;
    SS14[3][47] = 4'h0;
    SS14[4][47] = 4'h0;
    SS14[5][47] = 4'h0;
    SS14[6][47] = 4'h0;
    SS14[7][47] = 4'h0;
    SS14[8][47] = 4'h0;
    SS14[9][47] = 4'hD;
    SS14[10][47] = 4'hD;
    SS14[11][47] = 4'hD;
    SS14[12][47] = 4'h0;
    SS14[13][47] = 4'h0;
    SS14[14][47] = 4'h0;
    SS14[15][47] = 4'h0;
    SS14[16][47] = 4'h0;
    SS14[17][47] = 4'h0;
    SS14[18][47] = 4'h0;
    SS14[19][47] = 4'h0;
    SS14[20][47] = 4'h0;
    SS14[21][47] = 4'h0;
    SS14[22][47] = 4'h0;
    SS14[23][47] = 4'h0;
    SS14[24][47] = 4'h0;
    SS14[25][47] = 4'h0;
    SS14[26][47] = 4'h0;
    SS14[27][47] = 4'h0;
    SS14[28][47] = 4'h0;
    SS14[29][47] = 4'h0;
    SS14[30][47] = 4'h0;
    SS14[31][47] = 4'h0;
    SS14[32][47] = 4'h0;
    SS14[33][47] = 4'h0;
    SS14[34][47] = 4'h0;
    SS14[35][47] = 4'h0;
    SS14[36][47] = 4'hD;
    SS14[37][47] = 4'hD;
    SS14[38][47] = 4'hD;
    SS14[39][47] = 4'h0;
    SS14[40][47] = 4'h0;
    SS14[41][47] = 4'h0;
    SS14[42][47] = 4'h0;
    SS14[43][47] = 4'h0;
    SS14[44][47] = 4'h0;
    SS14[45][47] = 4'h0;
    SS14[46][47] = 4'h0;
    SS14[47][47] = 4'h0;
 
//SS 15
    SS15[0][0] = 4'h0;
    SS15[1][0] = 4'h0;
    SS15[2][0] = 4'h0;
    SS15[3][0] = 4'h0;
    SS15[4][0] = 4'h0;
    SS15[5][0] = 4'h0;
    SS15[6][0] = 4'h0;
    SS15[7][0] = 4'h0;
    SS15[8][0] = 4'h0;
    SS15[9][0] = 4'h0;
    SS15[10][0] = 4'h0;
    SS15[11][0] = 4'h0;
    SS15[12][0] = 4'h0;
    SS15[13][0] = 4'h0;
    SS15[14][0] = 4'h0;
    SS15[15][0] = 4'h0;
    SS15[16][0] = 4'h0;
    SS15[17][0] = 4'h0;
    SS15[18][0] = 4'h0;
    SS15[19][0] = 4'h0;
    SS15[20][0] = 4'h0;
    SS15[21][0] = 4'h0;
    SS15[22][0] = 4'h0;
    SS15[23][0] = 4'h0;
    SS15[24][0] = 4'h0;
    SS15[25][0] = 4'h0;
    SS15[26][0] = 4'h0;
    SS15[27][0] = 4'h0;
    SS15[28][0] = 4'h0;
    SS15[29][0] = 4'h0;
    SS15[30][0] = 4'h0;
    SS15[31][0] = 4'h0;
    SS15[32][0] = 4'h0;
    SS15[33][0] = 4'h0;
    SS15[34][0] = 4'h0;
    SS15[35][0] = 4'h0;
    SS15[36][0] = 4'h0;
    SS15[37][0] = 4'h0;
    SS15[38][0] = 4'h0;
    SS15[39][0] = 4'h0;
    SS15[40][0] = 4'h0;
    SS15[41][0] = 4'h0;
    SS15[42][0] = 4'h0;
    SS15[43][0] = 4'h0;
    SS15[44][0] = 4'h0;
    SS15[45][0] = 4'h0;
    SS15[46][0] = 4'h0;
    SS15[47][0] = 4'h0;
    SS15[0][1] = 4'h0;
    SS15[1][1] = 4'h0;
    SS15[2][1] = 4'h0;
    SS15[3][1] = 4'h0;
    SS15[4][1] = 4'h0;
    SS15[5][1] = 4'h0;
    SS15[6][1] = 4'h0;
    SS15[7][1] = 4'h0;
    SS15[8][1] = 4'h0;
    SS15[9][1] = 4'h0;
    SS15[10][1] = 4'h0;
    SS15[11][1] = 4'h0;
    SS15[12][1] = 4'h0;
    SS15[13][1] = 4'h0;
    SS15[14][1] = 4'h0;
    SS15[15][1] = 4'h0;
    SS15[16][1] = 4'h0;
    SS15[17][1] = 4'h0;
    SS15[18][1] = 4'h0;
    SS15[19][1] = 4'h0;
    SS15[20][1] = 4'h0;
    SS15[21][1] = 4'h0;
    SS15[22][1] = 4'h0;
    SS15[23][1] = 4'h0;
    SS15[24][1] = 4'h0;
    SS15[25][1] = 4'h0;
    SS15[26][1] = 4'h0;
    SS15[27][1] = 4'h0;
    SS15[28][1] = 4'h0;
    SS15[29][1] = 4'h0;
    SS15[30][1] = 4'hC;
    SS15[31][1] = 4'hC;
    SS15[32][1] = 4'h0;
    SS15[33][1] = 4'h0;
    SS15[34][1] = 4'h0;
    SS15[35][1] = 4'h0;
    SS15[36][1] = 4'h0;
    SS15[37][1] = 4'h0;
    SS15[38][1] = 4'h0;
    SS15[39][1] = 4'h0;
    SS15[40][1] = 4'h0;
    SS15[41][1] = 4'h0;
    SS15[42][1] = 4'h0;
    SS15[43][1] = 4'h0;
    SS15[44][1] = 4'h0;
    SS15[45][1] = 4'h0;
    SS15[46][1] = 4'h0;
    SS15[47][1] = 4'h0;
    SS15[0][2] = 4'h0;
    SS15[1][2] = 4'h0;
    SS15[2][2] = 4'h0;
    SS15[3][2] = 4'h0;
    SS15[4][2] = 4'h0;
    SS15[5][2] = 4'h0;
    SS15[6][2] = 4'h0;
    SS15[7][2] = 4'h0;
    SS15[8][2] = 4'h0;
    SS15[9][2] = 4'h0;
    SS15[10][2] = 4'h0;
    SS15[11][2] = 4'h0;
    SS15[12][2] = 4'h0;
    SS15[13][2] = 4'h0;
    SS15[14][2] = 4'h0;
    SS15[15][2] = 4'h0;
    SS15[16][2] = 4'h0;
    SS15[17][2] = 4'h0;
    SS15[18][2] = 4'h0;
    SS15[19][2] = 4'h0;
    SS15[20][2] = 4'h0;
    SS15[21][2] = 4'h0;
    SS15[22][2] = 4'h0;
    SS15[23][2] = 4'h0;
    SS15[24][2] = 4'h0;
    SS15[25][2] = 4'h0;
    SS15[26][2] = 4'h0;
    SS15[27][2] = 4'h0;
    SS15[28][2] = 4'h0;
    SS15[29][2] = 4'h0;
    SS15[30][2] = 4'hC;
    SS15[31][2] = 4'hC;
    SS15[32][2] = 4'hC;
    SS15[33][2] = 4'hC;
    SS15[34][2] = 4'h0;
    SS15[35][2] = 4'h0;
    SS15[36][2] = 4'h0;
    SS15[37][2] = 4'h0;
    SS15[38][2] = 4'h0;
    SS15[39][2] = 4'h0;
    SS15[40][2] = 4'h0;
    SS15[41][2] = 4'h0;
    SS15[42][2] = 4'h0;
    SS15[43][2] = 4'h0;
    SS15[44][2] = 4'h0;
    SS15[45][2] = 4'h0;
    SS15[46][2] = 4'h0;
    SS15[47][2] = 4'h0;
    SS15[0][3] = 4'h0;
    SS15[1][3] = 4'h0;
    SS15[2][3] = 4'h0;
    SS15[3][3] = 4'h0;
    SS15[4][3] = 4'h0;
    SS15[5][3] = 4'h0;
    SS15[6][3] = 4'h0;
    SS15[7][3] = 4'h0;
    SS15[8][3] = 4'h0;
    SS15[9][3] = 4'h0;
    SS15[10][3] = 4'h0;
    SS15[11][3] = 4'h0;
    SS15[12][3] = 4'h0;
    SS15[13][3] = 4'h0;
    SS15[14][3] = 4'h0;
    SS15[15][3] = 4'h0;
    SS15[16][3] = 4'h0;
    SS15[17][3] = 4'h0;
    SS15[18][3] = 4'h0;
    SS15[19][3] = 4'h0;
    SS15[20][3] = 4'h0;
    SS15[21][3] = 4'h0;
    SS15[22][3] = 4'h0;
    SS15[23][3] = 4'h0;
    SS15[24][3] = 4'h0;
    SS15[25][3] = 4'h0;
    SS15[26][3] = 4'h0;
    SS15[27][3] = 4'h0;
    SS15[28][3] = 4'h0;
    SS15[29][3] = 4'hC;
    SS15[30][3] = 4'hC;
    SS15[31][3] = 4'hC;
    SS15[32][3] = 4'hC;
    SS15[33][3] = 4'hC;
    SS15[34][3] = 4'hC;
    SS15[35][3] = 4'hC;
    SS15[36][3] = 4'h0;
    SS15[37][3] = 4'h0;
    SS15[38][3] = 4'h0;
    SS15[39][3] = 4'h0;
    SS15[40][3] = 4'h0;
    SS15[41][3] = 4'h0;
    SS15[42][3] = 4'h0;
    SS15[43][3] = 4'h0;
    SS15[44][3] = 4'h0;
    SS15[45][3] = 4'h0;
    SS15[46][3] = 4'h0;
    SS15[47][3] = 4'h0;
    SS15[0][4] = 4'h0;
    SS15[1][4] = 4'h0;
    SS15[2][4] = 4'h0;
    SS15[3][4] = 4'h0;
    SS15[4][4] = 4'h0;
    SS15[5][4] = 4'h0;
    SS15[6][4] = 4'h0;
    SS15[7][4] = 4'h0;
    SS15[8][4] = 4'h0;
    SS15[9][4] = 4'h0;
    SS15[10][4] = 4'h0;
    SS15[11][4] = 4'h0;
    SS15[12][4] = 4'h0;
    SS15[13][4] = 4'h0;
    SS15[14][4] = 4'h0;
    SS15[15][4] = 4'h0;
    SS15[16][4] = 4'h0;
    SS15[17][4] = 4'h0;
    SS15[18][4] = 4'h0;
    SS15[19][4] = 4'h0;
    SS15[20][4] = 4'h0;
    SS15[21][4] = 4'h0;
    SS15[22][4] = 4'h0;
    SS15[23][4] = 4'h0;
    SS15[24][4] = 4'h0;
    SS15[25][4] = 4'h0;
    SS15[26][4] = 4'h0;
    SS15[27][4] = 4'h0;
    SS15[28][4] = 4'h0;
    SS15[29][4] = 4'hC;
    SS15[30][4] = 4'hC;
    SS15[31][4] = 4'hC;
    SS15[32][4] = 4'hC;
    SS15[33][4] = 4'hC;
    SS15[34][4] = 4'hC;
    SS15[35][4] = 4'h0;
    SS15[36][4] = 4'h0;
    SS15[37][4] = 4'h0;
    SS15[38][4] = 4'h0;
    SS15[39][4] = 4'h0;
    SS15[40][4] = 4'h0;
    SS15[41][4] = 4'h0;
    SS15[42][4] = 4'h0;
    SS15[43][4] = 4'h0;
    SS15[44][4] = 4'h0;
    SS15[45][4] = 4'h0;
    SS15[46][4] = 4'h0;
    SS15[47][4] = 4'h0;
    SS15[0][5] = 4'h0;
    SS15[1][5] = 4'h0;
    SS15[2][5] = 4'h0;
    SS15[3][5] = 4'h0;
    SS15[4][5] = 4'h0;
    SS15[5][5] = 4'h0;
    SS15[6][5] = 4'h0;
    SS15[7][5] = 4'h0;
    SS15[8][5] = 4'h0;
    SS15[9][5] = 4'h0;
    SS15[10][5] = 4'h0;
    SS15[11][5] = 4'h0;
    SS15[12][5] = 4'h0;
    SS15[13][5] = 4'h0;
    SS15[14][5] = 4'h0;
    SS15[15][5] = 4'h0;
    SS15[16][5] = 4'h0;
    SS15[17][5] = 4'h0;
    SS15[18][5] = 4'h0;
    SS15[19][5] = 4'h0;
    SS15[20][5] = 4'h0;
    SS15[21][5] = 4'h0;
    SS15[22][5] = 4'h0;
    SS15[23][5] = 4'h0;
    SS15[24][5] = 4'h0;
    SS15[25][5] = 4'hD;
    SS15[26][5] = 4'h0;
    SS15[27][5] = 4'h0;
    SS15[28][5] = 4'hC;
    SS15[29][5] = 4'hC;
    SS15[30][5] = 4'hC;
    SS15[31][5] = 4'hC;
    SS15[32][5] = 4'hC;
    SS15[33][5] = 4'hC;
    SS15[34][5] = 4'hC;
    SS15[35][5] = 4'h0;
    SS15[36][5] = 4'h0;
    SS15[37][5] = 4'h0;
    SS15[38][5] = 4'h0;
    SS15[39][5] = 4'h0;
    SS15[40][5] = 4'h0;
    SS15[41][5] = 4'h0;
    SS15[42][5] = 4'h0;
    SS15[43][5] = 4'h0;
    SS15[44][5] = 4'h0;
    SS15[45][5] = 4'h0;
    SS15[46][5] = 4'h0;
    SS15[47][5] = 4'h0;
    SS15[0][6] = 4'h0;
    SS15[1][6] = 4'h0;
    SS15[2][6] = 4'h0;
    SS15[3][6] = 4'h0;
    SS15[4][6] = 4'h0;
    SS15[5][6] = 4'h0;
    SS15[6][6] = 4'h0;
    SS15[7][6] = 4'h0;
    SS15[8][6] = 4'h0;
    SS15[9][6] = 4'h0;
    SS15[10][6] = 4'h0;
    SS15[11][6] = 4'h0;
    SS15[12][6] = 4'h0;
    SS15[13][6] = 4'h0;
    SS15[14][6] = 4'h0;
    SS15[15][6] = 4'h0;
    SS15[16][6] = 4'h0;
    SS15[17][6] = 4'h0;
    SS15[18][6] = 4'h0;
    SS15[19][6] = 4'h0;
    SS15[20][6] = 4'h0;
    SS15[21][6] = 4'h0;
    SS15[22][6] = 4'h0;
    SS15[23][6] = 4'h0;
    SS15[24][6] = 4'h0;
    SS15[25][6] = 4'hD;
    SS15[26][6] = 4'hD;
    SS15[27][6] = 4'hD;
    SS15[28][6] = 4'hC;
    SS15[29][6] = 4'hC;
    SS15[30][6] = 4'hC;
    SS15[31][6] = 4'hC;
    SS15[32][6] = 4'hC;
    SS15[33][6] = 4'hC;
    SS15[34][6] = 4'h0;
    SS15[35][6] = 4'h0;
    SS15[36][6] = 4'h0;
    SS15[37][6] = 4'h0;
    SS15[38][6] = 4'h0;
    SS15[39][6] = 4'h0;
    SS15[40][6] = 4'h0;
    SS15[41][6] = 4'h0;
    SS15[42][6] = 4'h0;
    SS15[43][6] = 4'h0;
    SS15[44][6] = 4'h0;
    SS15[45][6] = 4'h0;
    SS15[46][6] = 4'h0;
    SS15[47][6] = 4'h0;
    SS15[0][7] = 4'h0;
    SS15[1][7] = 4'h0;
    SS15[2][7] = 4'h0;
    SS15[3][7] = 4'h0;
    SS15[4][7] = 4'h0;
    SS15[5][7] = 4'h0;
    SS15[6][7] = 4'h0;
    SS15[7][7] = 4'h0;
    SS15[8][7] = 4'h0;
    SS15[9][7] = 4'h0;
    SS15[10][7] = 4'h0;
    SS15[11][7] = 4'h0;
    SS15[12][7] = 4'h0;
    SS15[13][7] = 4'h0;
    SS15[14][7] = 4'h0;
    SS15[15][7] = 4'h0;
    SS15[16][7] = 4'h0;
    SS15[17][7] = 4'h0;
    SS15[18][7] = 4'h0;
    SS15[19][7] = 4'h0;
    SS15[20][7] = 4'h0;
    SS15[21][7] = 4'h0;
    SS15[22][7] = 4'h0;
    SS15[23][7] = 4'h0;
    SS15[24][7] = 4'hD;
    SS15[25][7] = 4'hD;
    SS15[26][7] = 4'hD;
    SS15[27][7] = 4'hD;
    SS15[28][7] = 4'hC;
    SS15[29][7] = 4'hC;
    SS15[30][7] = 4'hC;
    SS15[31][7] = 4'hC;
    SS15[32][7] = 4'hC;
    SS15[33][7] = 4'hC;
    SS15[34][7] = 4'h0;
    SS15[35][7] = 4'h0;
    SS15[36][7] = 4'h0;
    SS15[37][7] = 4'h0;
    SS15[38][7] = 4'h0;
    SS15[39][7] = 4'h0;
    SS15[40][7] = 4'h0;
    SS15[41][7] = 4'h0;
    SS15[42][7] = 4'h0;
    SS15[43][7] = 4'h0;
    SS15[44][7] = 4'h0;
    SS15[45][7] = 4'h0;
    SS15[46][7] = 4'h0;
    SS15[47][7] = 4'h0;
    SS15[0][8] = 4'h0;
    SS15[1][8] = 4'h0;
    SS15[2][8] = 4'h0;
    SS15[3][8] = 4'h0;
    SS15[4][8] = 4'h0;
    SS15[5][8] = 4'h0;
    SS15[6][8] = 4'h0;
    SS15[7][8] = 4'h0;
    SS15[8][8] = 4'h0;
    SS15[9][8] = 4'h0;
    SS15[10][8] = 4'h0;
    SS15[11][8] = 4'h0;
    SS15[12][8] = 4'h0;
    SS15[13][8] = 4'h0;
    SS15[14][8] = 4'h0;
    SS15[15][8] = 4'h0;
    SS15[16][8] = 4'h0;
    SS15[17][8] = 4'h0;
    SS15[18][8] = 4'h0;
    SS15[19][8] = 4'h0;
    SS15[20][8] = 4'h0;
    SS15[21][8] = 4'h0;
    SS15[22][8] = 4'h0;
    SS15[23][8] = 4'h0;
    SS15[24][8] = 4'hD;
    SS15[25][8] = 4'hD;
    SS15[26][8] = 4'hD;
    SS15[27][8] = 4'hC;
    SS15[28][8] = 4'hC;
    SS15[29][8] = 4'hC;
    SS15[30][8] = 4'hC;
    SS15[31][8] = 4'hC;
    SS15[32][8] = 4'hC;
    SS15[33][8] = 4'hC;
    SS15[34][8] = 4'h0;
    SS15[35][8] = 4'h0;
    SS15[36][8] = 4'h0;
    SS15[37][8] = 4'h0;
    SS15[38][8] = 4'h0;
    SS15[39][8] = 4'h0;
    SS15[40][8] = 4'h0;
    SS15[41][8] = 4'h0;
    SS15[42][8] = 4'h0;
    SS15[43][8] = 4'h0;
    SS15[44][8] = 4'h0;
    SS15[45][8] = 4'h0;
    SS15[46][8] = 4'h0;
    SS15[47][8] = 4'h0;
    SS15[0][9] = 4'h0;
    SS15[1][9] = 4'h0;
    SS15[2][9] = 4'h0;
    SS15[3][9] = 4'h0;
    SS15[4][9] = 4'h0;
    SS15[5][9] = 4'h0;
    SS15[6][9] = 4'h0;
    SS15[7][9] = 4'h0;
    SS15[8][9] = 4'h0;
    SS15[9][9] = 4'h0;
    SS15[10][9] = 4'h0;
    SS15[11][9] = 4'h0;
    SS15[12][9] = 4'h0;
    SS15[13][9] = 4'h0;
    SS15[14][9] = 4'h0;
    SS15[15][9] = 4'h0;
    SS15[16][9] = 4'h0;
    SS15[17][9] = 4'h0;
    SS15[18][9] = 4'h0;
    SS15[19][9] = 4'h0;
    SS15[20][9] = 4'h0;
    SS15[21][9] = 4'h0;
    SS15[22][9] = 4'h0;
    SS15[23][9] = 4'h0;
    SS15[24][9] = 4'hD;
    SS15[25][9] = 4'hD;
    SS15[26][9] = 4'hD;
    SS15[27][9] = 4'hC;
    SS15[28][9] = 4'hC;
    SS15[29][9] = 4'hC;
    SS15[30][9] = 4'hC;
    SS15[31][9] = 4'hC;
    SS15[32][9] = 4'hC;
    SS15[33][9] = 4'hD;
    SS15[34][9] = 4'hD;
    SS15[35][9] = 4'hF;
    SS15[36][9] = 4'h0;
    SS15[37][9] = 4'h0;
    SS15[38][9] = 4'h0;
    SS15[39][9] = 4'h0;
    SS15[40][9] = 4'h0;
    SS15[41][9] = 4'h0;
    SS15[42][9] = 4'h0;
    SS15[43][9] = 4'h0;
    SS15[44][9] = 4'h0;
    SS15[45][9] = 4'h0;
    SS15[46][9] = 4'h0;
    SS15[47][9] = 4'h0;
    SS15[0][10] = 4'h0;
    SS15[1][10] = 4'h0;
    SS15[2][10] = 4'h0;
    SS15[3][10] = 4'h0;
    SS15[4][10] = 4'h0;
    SS15[5][10] = 4'h0;
    SS15[6][10] = 4'h0;
    SS15[7][10] = 4'h0;
    SS15[8][10] = 4'h0;
    SS15[9][10] = 4'h0;
    SS15[10][10] = 4'h0;
    SS15[11][10] = 4'h0;
    SS15[12][10] = 4'h0;
    SS15[13][10] = 4'h0;
    SS15[14][10] = 4'h0;
    SS15[15][10] = 4'h0;
    SS15[16][10] = 4'h0;
    SS15[17][10] = 4'h0;
    SS15[18][10] = 4'h0;
    SS15[19][10] = 4'h0;
    SS15[20][10] = 4'h0;
    SS15[21][10] = 4'h0;
    SS15[22][10] = 4'h0;
    SS15[23][10] = 4'hD;
    SS15[24][10] = 4'hD;
    SS15[25][10] = 4'hD;
    SS15[26][10] = 4'hC;
    SS15[27][10] = 4'hC;
    SS15[28][10] = 4'hC;
    SS15[29][10] = 4'hC;
    SS15[30][10] = 4'hC;
    SS15[31][10] = 4'hC;
    SS15[32][10] = 4'hC;
    SS15[33][10] = 4'hD;
    SS15[34][10] = 4'hD;
    SS15[35][10] = 4'hD;
    SS15[36][10] = 4'h0;
    SS15[37][10] = 4'h0;
    SS15[38][10] = 4'h0;
    SS15[39][10] = 4'h0;
    SS15[40][10] = 4'h0;
    SS15[41][10] = 4'h0;
    SS15[42][10] = 4'h0;
    SS15[43][10] = 4'h0;
    SS15[44][10] = 4'h0;
    SS15[45][10] = 4'h0;
    SS15[46][10] = 4'h0;
    SS15[47][10] = 4'h0;
    SS15[0][11] = 4'h0;
    SS15[1][11] = 4'h0;
    SS15[2][11] = 4'h0;
    SS15[3][11] = 4'h0;
    SS15[4][11] = 4'h0;
    SS15[5][11] = 4'h0;
    SS15[6][11] = 4'h0;
    SS15[7][11] = 4'h0;
    SS15[8][11] = 4'h0;
    SS15[9][11] = 4'h0;
    SS15[10][11] = 4'h0;
    SS15[11][11] = 4'h0;
    SS15[12][11] = 4'h0;
    SS15[13][11] = 4'h0;
    SS15[14][11] = 4'h0;
    SS15[15][11] = 4'h0;
    SS15[16][11] = 4'h0;
    SS15[17][11] = 4'h0;
    SS15[18][11] = 4'h0;
    SS15[19][11] = 4'h0;
    SS15[20][11] = 4'h0;
    SS15[21][11] = 4'h0;
    SS15[22][11] = 4'h0;
    SS15[23][11] = 4'hD;
    SS15[24][11] = 4'hD;
    SS15[25][11] = 4'hD;
    SS15[26][11] = 4'hC;
    SS15[27][11] = 4'hC;
    SS15[28][11] = 4'hC;
    SS15[29][11] = 4'hC;
    SS15[30][11] = 4'hC;
    SS15[31][11] = 4'hC;
    SS15[32][11] = 4'hD;
    SS15[33][11] = 4'hD;
    SS15[34][11] = 4'hD;
    SS15[35][11] = 4'hD;
    SS15[36][11] = 4'h0;
    SS15[37][11] = 4'h0;
    SS15[38][11] = 4'h0;
    SS15[39][11] = 4'h0;
    SS15[40][11] = 4'h0;
    SS15[41][11] = 4'h0;
    SS15[42][11] = 4'h0;
    SS15[43][11] = 4'h0;
    SS15[44][11] = 4'h0;
    SS15[45][11] = 4'h0;
    SS15[46][11] = 4'h0;
    SS15[47][11] = 4'h0;
    SS15[0][12] = 4'h0;
    SS15[1][12] = 4'h0;
    SS15[2][12] = 4'h0;
    SS15[3][12] = 4'h0;
    SS15[4][12] = 4'h0;
    SS15[5][12] = 4'h0;
    SS15[6][12] = 4'h0;
    SS15[7][12] = 4'h0;
    SS15[8][12] = 4'h0;
    SS15[9][12] = 4'h0;
    SS15[10][12] = 4'h0;
    SS15[11][12] = 4'h0;
    SS15[12][12] = 4'h0;
    SS15[13][12] = 4'h0;
    SS15[14][12] = 4'h0;
    SS15[15][12] = 4'h0;
    SS15[16][12] = 4'h0;
    SS15[17][12] = 4'h0;
    SS15[18][12] = 4'h0;
    SS15[19][12] = 4'h0;
    SS15[20][12] = 4'h0;
    SS15[21][12] = 4'h0;
    SS15[22][12] = 4'hD;
    SS15[23][12] = 4'hD;
    SS15[24][12] = 4'hD;
    SS15[25][12] = 4'hD;
    SS15[26][12] = 4'hC;
    SS15[27][12] = 4'hC;
    SS15[28][12] = 4'hC;
    SS15[29][12] = 4'hC;
    SS15[30][12] = 4'hC;
    SS15[31][12] = 4'hC;
    SS15[32][12] = 4'hD;
    SS15[33][12] = 4'hD;
    SS15[34][12] = 4'hD;
    SS15[35][12] = 4'h0;
    SS15[36][12] = 4'h0;
    SS15[37][12] = 4'h0;
    SS15[38][12] = 4'h0;
    SS15[39][12] = 4'h0;
    SS15[40][12] = 4'h0;
    SS15[41][12] = 4'h0;
    SS15[42][12] = 4'h0;
    SS15[43][12] = 4'h0;
    SS15[44][12] = 4'h0;
    SS15[45][12] = 4'h0;
    SS15[46][12] = 4'h0;
    SS15[47][12] = 4'h0;
    SS15[0][13] = 4'h0;
    SS15[1][13] = 4'h0;
    SS15[2][13] = 4'h0;
    SS15[3][13] = 4'h0;
    SS15[4][13] = 4'h0;
    SS15[5][13] = 4'h0;
    SS15[6][13] = 4'h0;
    SS15[7][13] = 4'h0;
    SS15[8][13] = 4'h0;
    SS15[9][13] = 4'h0;
    SS15[10][13] = 4'h0;
    SS15[11][13] = 4'h0;
    SS15[12][13] = 4'h0;
    SS15[13][13] = 4'h0;
    SS15[14][13] = 4'h0;
    SS15[15][13] = 4'h0;
    SS15[16][13] = 4'h0;
    SS15[17][13] = 4'h0;
    SS15[18][13] = 4'h0;
    SS15[19][13] = 4'h0;
    SS15[20][13] = 4'h0;
    SS15[21][13] = 4'h0;
    SS15[22][13] = 4'hD;
    SS15[23][13] = 4'hD;
    SS15[24][13] = 4'hD;
    SS15[25][13] = 4'hC;
    SS15[26][13] = 4'hC;
    SS15[27][13] = 4'hC;
    SS15[28][13] = 4'hC;
    SS15[29][13] = 4'hC;
    SS15[30][13] = 4'hC;
    SS15[31][13] = 4'hC;
    SS15[32][13] = 4'hD;
    SS15[33][13] = 4'hD;
    SS15[34][13] = 4'hD;
    SS15[35][13] = 4'h0;
    SS15[36][13] = 4'h0;
    SS15[37][13] = 4'h0;
    SS15[38][13] = 4'h0;
    SS15[39][13] = 4'h0;
    SS15[40][13] = 4'h0;
    SS15[41][13] = 4'h0;
    SS15[42][13] = 4'h0;
    SS15[43][13] = 4'h0;
    SS15[44][13] = 4'h0;
    SS15[45][13] = 4'h0;
    SS15[46][13] = 4'h0;
    SS15[47][13] = 4'h0;
    SS15[0][14] = 4'h0;
    SS15[1][14] = 4'h0;
    SS15[2][14] = 4'h0;
    SS15[3][14] = 4'h0;
    SS15[4][14] = 4'h0;
    SS15[5][14] = 4'h0;
    SS15[6][14] = 4'h0;
    SS15[7][14] = 4'h0;
    SS15[8][14] = 4'h0;
    SS15[9][14] = 4'h0;
    SS15[10][14] = 4'h0;
    SS15[11][14] = 4'h0;
    SS15[12][14] = 4'h0;
    SS15[13][14] = 4'h0;
    SS15[14][14] = 4'h0;
    SS15[15][14] = 4'h3;
    SS15[16][14] = 4'h3;
    SS15[17][14] = 4'h0;
    SS15[18][14] = 4'h0;
    SS15[19][14] = 4'h0;
    SS15[20][14] = 4'h0;
    SS15[21][14] = 4'hE;
    SS15[22][14] = 4'hC;
    SS15[23][14] = 4'hC;
    SS15[24][14] = 4'hD;
    SS15[25][14] = 4'hC;
    SS15[26][14] = 4'hC;
    SS15[27][14] = 4'hC;
    SS15[28][14] = 4'hC;
    SS15[29][14] = 4'hC;
    SS15[30][14] = 4'hC;
    SS15[31][14] = 4'hD;
    SS15[32][14] = 4'hD;
    SS15[33][14] = 4'hD;
    SS15[34][14] = 4'h0;
    SS15[35][14] = 4'h0;
    SS15[36][14] = 4'h0;
    SS15[37][14] = 4'h0;
    SS15[38][14] = 4'h0;
    SS15[39][14] = 4'h0;
    SS15[40][14] = 4'h0;
    SS15[41][14] = 4'h0;
    SS15[42][14] = 4'h0;
    SS15[43][14] = 4'h0;
    SS15[44][14] = 4'h0;
    SS15[45][14] = 4'h0;
    SS15[46][14] = 4'h0;
    SS15[47][14] = 4'h0;
    SS15[0][15] = 4'h0;
    SS15[1][15] = 4'h0;
    SS15[2][15] = 4'h0;
    SS15[3][15] = 4'h0;
    SS15[4][15] = 4'h0;
    SS15[5][15] = 4'h0;
    SS15[6][15] = 4'h0;
    SS15[7][15] = 4'h0;
    SS15[8][15] = 4'h0;
    SS15[9][15] = 4'h0;
    SS15[10][15] = 4'h0;
    SS15[11][15] = 4'h0;
    SS15[12][15] = 4'h0;
    SS15[13][15] = 4'h0;
    SS15[14][15] = 4'h0;
    SS15[15][15] = 4'h3;
    SS15[16][15] = 4'h3;
    SS15[17][15] = 4'h3;
    SS15[18][15] = 4'hD;
    SS15[19][15] = 4'h0;
    SS15[20][15] = 4'h0;
    SS15[21][15] = 4'hC;
    SS15[22][15] = 4'hC;
    SS15[23][15] = 4'hC;
    SS15[24][15] = 4'hC;
    SS15[25][15] = 4'hC;
    SS15[26][15] = 4'hC;
    SS15[27][15] = 4'hC;
    SS15[28][15] = 4'hC;
    SS15[29][15] = 4'hC;
    SS15[30][15] = 4'hC;
    SS15[31][15] = 4'hD;
    SS15[32][15] = 4'hD;
    SS15[33][15] = 4'hD;
    SS15[34][15] = 4'h0;
    SS15[35][15] = 4'h0;
    SS15[36][15] = 4'h0;
    SS15[37][15] = 4'h0;
    SS15[38][15] = 4'h0;
    SS15[39][15] = 4'h0;
    SS15[40][15] = 4'h0;
    SS15[41][15] = 4'h0;
    SS15[42][15] = 4'h0;
    SS15[43][15] = 4'h0;
    SS15[44][15] = 4'h0;
    SS15[45][15] = 4'h0;
    SS15[46][15] = 4'h0;
    SS15[47][15] = 4'h0;
    SS15[0][16] = 4'h0;
    SS15[1][16] = 4'h0;
    SS15[2][16] = 4'h0;
    SS15[3][16] = 4'h0;
    SS15[4][16] = 4'h0;
    SS15[5][16] = 4'h0;
    SS15[6][16] = 4'h0;
    SS15[7][16] = 4'h0;
    SS15[8][16] = 4'h0;
    SS15[9][16] = 4'h0;
    SS15[10][16] = 4'h0;
    SS15[11][16] = 4'h0;
    SS15[12][16] = 4'h0;
    SS15[13][16] = 4'h0;
    SS15[14][16] = 4'h3;
    SS15[15][16] = 4'h3;
    SS15[16][16] = 4'h3;
    SS15[17][16] = 4'hD;
    SS15[18][16] = 4'hD;
    SS15[19][16] = 4'hD;
    SS15[20][16] = 4'hD;
    SS15[21][16] = 4'hC;
    SS15[22][16] = 4'hC;
    SS15[23][16] = 4'hC;
    SS15[24][16] = 4'hC;
    SS15[25][16] = 4'hC;
    SS15[26][16] = 4'hC;
    SS15[27][16] = 4'hC;
    SS15[28][16] = 4'hC;
    SS15[29][16] = 4'hC;
    SS15[30][16] = 4'hD;
    SS15[31][16] = 4'hD;
    SS15[32][16] = 4'hD;
    SS15[33][16] = 4'hD;
    SS15[34][16] = 4'h0;
    SS15[35][16] = 4'h0;
    SS15[36][16] = 4'h0;
    SS15[37][16] = 4'h0;
    SS15[38][16] = 4'h0;
    SS15[39][16] = 4'h0;
    SS15[40][16] = 4'h0;
    SS15[41][16] = 4'h0;
    SS15[42][16] = 4'h0;
    SS15[43][16] = 4'h0;
    SS15[44][16] = 4'h0;
    SS15[45][16] = 4'h0;
    SS15[46][16] = 4'h0;
    SS15[47][16] = 4'h0;
    SS15[0][17] = 4'h0;
    SS15[1][17] = 4'h0;
    SS15[2][17] = 4'h0;
    SS15[3][17] = 4'h0;
    SS15[4][17] = 4'h0;
    SS15[5][17] = 4'h0;
    SS15[6][17] = 4'h0;
    SS15[7][17] = 4'h3;
    SS15[8][17] = 4'h0;
    SS15[9][17] = 4'h0;
    SS15[10][17] = 4'h0;
    SS15[11][17] = 4'h0;
    SS15[12][17] = 4'h0;
    SS15[13][17] = 4'h0;
    SS15[14][17] = 4'hD;
    SS15[15][17] = 4'hD;
    SS15[16][17] = 4'h3;
    SS15[17][17] = 4'hD;
    SS15[18][17] = 4'hD;
    SS15[19][17] = 4'hD;
    SS15[20][17] = 4'hD;
    SS15[21][17] = 4'hD;
    SS15[22][17] = 4'hD;
    SS15[23][17] = 4'hA;
    SS15[24][17] = 4'hC;
    SS15[25][17] = 4'hC;
    SS15[26][17] = 4'hC;
    SS15[27][17] = 4'hC;
    SS15[28][17] = 4'hC;
    SS15[29][17] = 4'hC;
    SS15[30][17] = 4'hC;
    SS15[31][17] = 4'hC;
    SS15[32][17] = 4'hD;
    SS15[33][17] = 4'h0;
    SS15[34][17] = 4'h0;
    SS15[35][17] = 4'h0;
    SS15[36][17] = 4'h0;
    SS15[37][17] = 4'h0;
    SS15[38][17] = 4'h0;
    SS15[39][17] = 4'h0;
    SS15[40][17] = 4'h0;
    SS15[41][17] = 4'h0;
    SS15[42][17] = 4'h0;
    SS15[43][17] = 4'h0;
    SS15[44][17] = 4'h0;
    SS15[45][17] = 4'h0;
    SS15[46][17] = 4'h0;
    SS15[47][17] = 4'h0;
    SS15[0][18] = 4'h0;
    SS15[1][18] = 4'h0;
    SS15[2][18] = 4'h0;
    SS15[3][18] = 4'h0;
    SS15[4][18] = 4'h0;
    SS15[5][18] = 4'h0;
    SS15[6][18] = 4'h0;
    SS15[7][18] = 4'h3;
    SS15[8][18] = 4'h3;
    SS15[9][18] = 4'h3;
    SS15[10][18] = 4'hD;
    SS15[11][18] = 4'h0;
    SS15[12][18] = 4'h0;
    SS15[13][18] = 4'hD;
    SS15[14][18] = 4'hD;
    SS15[15][18] = 4'hD;
    SS15[16][18] = 4'hD;
    SS15[17][18] = 4'hD;
    SS15[18][18] = 4'hD;
    SS15[19][18] = 4'hD;
    SS15[20][18] = 4'hD;
    SS15[21][18] = 4'hD;
    SS15[22][18] = 4'hD;
    SS15[23][18] = 4'hA;
    SS15[24][18] = 4'hA;
    SS15[25][18] = 4'hA;
    SS15[26][18] = 4'hC;
    SS15[27][18] = 4'hC;
    SS15[28][18] = 4'hC;
    SS15[29][18] = 4'hC;
    SS15[30][18] = 4'hC;
    SS15[31][18] = 4'hC;
    SS15[32][18] = 4'hC;
    SS15[33][18] = 4'h0;
    SS15[34][18] = 4'h0;
    SS15[35][18] = 4'h0;
    SS15[36][18] = 4'h0;
    SS15[37][18] = 4'h0;
    SS15[38][18] = 4'h0;
    SS15[39][18] = 4'h0;
    SS15[40][18] = 4'h0;
    SS15[41][18] = 4'h0;
    SS15[42][18] = 4'h0;
    SS15[43][18] = 4'h0;
    SS15[44][18] = 4'h0;
    SS15[45][18] = 4'h0;
    SS15[46][18] = 4'h0;
    SS15[47][18] = 4'h0;
    SS15[0][19] = 4'h0;
    SS15[1][19] = 4'h0;
    SS15[2][19] = 4'h0;
    SS15[3][19] = 4'hD;
    SS15[4][19] = 4'hD;
    SS15[5][19] = 4'h0;
    SS15[6][19] = 4'h0;
    SS15[7][19] = 4'h3;
    SS15[8][19] = 4'h3;
    SS15[9][19] = 4'h3;
    SS15[10][19] = 4'hD;
    SS15[11][19] = 4'hD;
    SS15[12][19] = 4'hD;
    SS15[13][19] = 4'hD;
    SS15[14][19] = 4'hD;
    SS15[15][19] = 4'hD;
    SS15[16][19] = 4'hD;
    SS15[17][19] = 4'hD;
    SS15[18][19] = 4'hD;
    SS15[19][19] = 4'hC;
    SS15[20][19] = 4'hC;
    SS15[21][19] = 4'hD;
    SS15[22][19] = 4'hD;
    SS15[23][19] = 4'hA;
    SS15[24][19] = 4'hA;
    SS15[25][19] = 4'hA;
    SS15[26][19] = 4'hA;
    SS15[27][19] = 4'hA;
    SS15[28][19] = 4'hA;
    SS15[29][19] = 4'hC;
    SS15[30][19] = 4'hC;
    SS15[31][19] = 4'hC;
    SS15[32][19] = 4'h0;
    SS15[33][19] = 4'h0;
    SS15[34][19] = 4'h0;
    SS15[35][19] = 4'h0;
    SS15[36][19] = 4'h0;
    SS15[37][19] = 4'h0;
    SS15[38][19] = 4'h0;
    SS15[39][19] = 4'h0;
    SS15[40][19] = 4'h0;
    SS15[41][19] = 4'h0;
    SS15[42][19] = 4'h0;
    SS15[43][19] = 4'h0;
    SS15[44][19] = 4'h0;
    SS15[45][19] = 4'h0;
    SS15[46][19] = 4'h0;
    SS15[47][19] = 4'h0;
    SS15[0][20] = 4'h0;
    SS15[1][20] = 4'h0;
    SS15[2][20] = 4'h0;
    SS15[3][20] = 4'hD;
    SS15[4][20] = 4'hD;
    SS15[5][20] = 4'hD;
    SS15[6][20] = 4'hD;
    SS15[7][20] = 4'hD;
    SS15[8][20] = 4'h3;
    SS15[9][20] = 4'hD;
    SS15[10][20] = 4'hD;
    SS15[11][20] = 4'hD;
    SS15[12][20] = 4'hD;
    SS15[13][20] = 4'hD;
    SS15[14][20] = 4'hD;
    SS15[15][20] = 4'hD;
    SS15[16][20] = 4'hD;
    SS15[17][20] = 4'hD;
    SS15[18][20] = 4'hD;
    SS15[19][20] = 4'hC;
    SS15[20][20] = 4'hC;
    SS15[21][20] = 4'hC;
    SS15[22][20] = 4'hD;
    SS15[23][20] = 4'hA;
    SS15[24][20] = 4'hA;
    SS15[25][20] = 4'hA;
    SS15[26][20] = 4'hA;
    SS15[27][20] = 4'hA;
    SS15[28][20] = 4'hA;
    SS15[29][20] = 4'hD;
    SS15[30][20] = 4'hD;
    SS15[31][20] = 4'hC;
    SS15[32][20] = 4'h0;
    SS15[33][20] = 4'h0;
    SS15[34][20] = 4'h0;
    SS15[35][20] = 4'h0;
    SS15[36][20] = 4'h0;
    SS15[37][20] = 4'h0;
    SS15[38][20] = 4'h0;
    SS15[39][20] = 4'h0;
    SS15[40][20] = 4'h0;
    SS15[41][20] = 4'h0;
    SS15[42][20] = 4'h0;
    SS15[43][20] = 4'h0;
    SS15[44][20] = 4'h0;
    SS15[45][20] = 4'h0;
    SS15[46][20] = 4'h0;
    SS15[47][20] = 4'h0;
    SS15[0][21] = 4'hD;
    SS15[1][21] = 4'hD;
    SS15[2][21] = 4'hE;
    SS15[3][21] = 4'hD;
    SS15[4][21] = 4'hD;
    SS15[5][21] = 4'hD;
    SS15[6][21] = 4'hD;
    SS15[7][21] = 4'hD;
    SS15[8][21] = 4'hD;
    SS15[9][21] = 4'hE;
    SS15[10][21] = 4'hD;
    SS15[11][21] = 4'hD;
    SS15[12][21] = 4'hD;
    SS15[13][21] = 4'hD;
    SS15[14][21] = 4'hD;
    SS15[15][21] = 4'hE;
    SS15[16][21] = 4'hE;
    SS15[17][21] = 4'hE;
    SS15[18][21] = 4'hD;
    SS15[19][21] = 4'hC;
    SS15[20][21] = 4'hC;
    SS15[21][21] = 4'hC;
    SS15[22][21] = 4'hD;
    SS15[23][21] = 4'hD;
    SS15[24][21] = 4'hD;
    SS15[25][21] = 4'hD;
    SS15[26][21] = 4'hA;
    SS15[27][21] = 4'hA;
    SS15[28][21] = 4'hD;
    SS15[29][21] = 4'hD;
    SS15[30][21] = 4'hD;
    SS15[31][21] = 4'hD;
    SS15[32][21] = 4'hD;
    SS15[33][21] = 4'hF;
    SS15[34][21] = 4'h0;
    SS15[35][21] = 4'h0;
    SS15[36][21] = 4'h0;
    SS15[37][21] = 4'h0;
    SS15[38][21] = 4'h0;
    SS15[39][21] = 4'h0;
    SS15[40][21] = 4'h0;
    SS15[41][21] = 4'h0;
    SS15[42][21] = 4'h0;
    SS15[43][21] = 4'h0;
    SS15[44][21] = 4'h0;
    SS15[45][21] = 4'h0;
    SS15[46][21] = 4'h0;
    SS15[47][21] = 4'h0;
    SS15[0][22] = 4'hD;
    SS15[1][22] = 4'hD;
    SS15[2][22] = 4'hD;
    SS15[3][22] = 4'hD;
    SS15[4][22] = 4'hD;
    SS15[5][22] = 4'hD;
    SS15[6][22] = 4'hD;
    SS15[7][22] = 4'hD;
    SS15[8][22] = 4'hD;
    SS15[9][22] = 4'hE;
    SS15[10][22] = 4'hE;
    SS15[11][22] = 4'hE;
    SS15[12][22] = 4'hE;
    SS15[13][22] = 4'hD;
    SS15[14][22] = 4'hD;
    SS15[15][22] = 4'hE;
    SS15[16][22] = 4'hE;
    SS15[17][22] = 4'hE;
    SS15[18][22] = 4'hC;
    SS15[19][22] = 4'hC;
    SS15[20][22] = 4'hC;
    SS15[21][22] = 4'hD;
    SS15[22][22] = 4'hD;
    SS15[23][22] = 4'hD;
    SS15[24][22] = 4'hD;
    SS15[25][22] = 4'hD;
    SS15[26][22] = 4'hD;
    SS15[27][22] = 4'hD;
    SS15[28][22] = 4'hD;
    SS15[29][22] = 4'hD;
    SS15[30][22] = 4'hD;
    SS15[31][22] = 4'hD;
    SS15[32][22] = 4'hD;
    SS15[33][22] = 4'hD;
    SS15[34][22] = 4'h3;
    SS15[35][22] = 4'h3;
    SS15[36][22] = 4'h0;
    SS15[37][22] = 4'h0;
    SS15[38][22] = 4'h0;
    SS15[39][22] = 4'h0;
    SS15[40][22] = 4'h0;
    SS15[41][22] = 4'h0;
    SS15[42][22] = 4'h0;
    SS15[43][22] = 4'h0;
    SS15[44][22] = 4'h0;
    SS15[45][22] = 4'h0;
    SS15[46][22] = 4'h0;
    SS15[47][22] = 4'h0;
    SS15[0][23] = 4'hD;
    SS15[1][23] = 4'hD;
    SS15[2][23] = 4'hD;
    SS15[3][23] = 4'hD;
    SS15[4][23] = 4'hD;
    SS15[5][23] = 4'hE;
    SS15[6][23] = 4'hE;
    SS15[7][23] = 4'hD;
    SS15[8][23] = 4'hE;
    SS15[9][23] = 4'hE;
    SS15[10][23] = 4'hE;
    SS15[11][23] = 4'hE;
    SS15[12][23] = 4'hE;
    SS15[13][23] = 4'hE;
    SS15[14][23] = 4'hE;
    SS15[15][23] = 4'hE;
    SS15[16][23] = 4'hE;
    SS15[17][23] = 4'hE;
    SS15[18][23] = 4'hC;
    SS15[19][23] = 4'hC;
    SS15[20][23] = 4'hC;
    SS15[21][23] = 4'hC;
    SS15[22][23] = 4'hC;
    SS15[23][23] = 4'hD;
    SS15[24][23] = 4'hD;
    SS15[25][23] = 4'hD;
    SS15[26][23] = 4'hD;
    SS15[27][23] = 4'hC;
    SS15[28][23] = 4'hC;
    SS15[29][23] = 4'hC;
    SS15[30][23] = 4'hC;
    SS15[31][23] = 4'hD;
    SS15[32][23] = 4'hD;
    SS15[33][23] = 4'hD;
    SS15[34][23] = 4'h3;
    SS15[35][23] = 4'h3;
    SS15[36][23] = 4'h3;
    SS15[37][23] = 4'h0;
    SS15[38][23] = 4'h0;
    SS15[39][23] = 4'h0;
    SS15[40][23] = 4'h0;
    SS15[41][23] = 4'h0;
    SS15[42][23] = 4'h0;
    SS15[43][23] = 4'h0;
    SS15[44][23] = 4'h0;
    SS15[45][23] = 4'h0;
    SS15[46][23] = 4'h0;
    SS15[47][23] = 4'h0;
    SS15[0][24] = 4'h0;
    SS15[1][24] = 4'h0;
    SS15[2][24] = 4'hD;
    SS15[3][24] = 4'hD;
    SS15[4][24] = 4'hD;
    SS15[5][24] = 4'hE;
    SS15[6][24] = 4'hE;
    SS15[7][24] = 4'hE;
    SS15[8][24] = 4'hE;
    SS15[9][24] = 4'hE;
    SS15[10][24] = 4'hE;
    SS15[11][24] = 4'hE;
    SS15[12][24] = 4'hE;
    SS15[13][24] = 4'hE;
    SS15[14][24] = 4'hC;
    SS15[15][24] = 4'hC;
    SS15[16][24] = 4'hC;
    SS15[17][24] = 4'hC;
    SS15[18][24] = 4'hC;
    SS15[19][24] = 4'hC;
    SS15[20][24] = 4'hC;
    SS15[21][24] = 4'hC;
    SS15[22][24] = 4'hC;
    SS15[23][24] = 4'hC;
    SS15[24][24] = 4'hC;
    SS15[25][24] = 4'hD;
    SS15[26][24] = 4'hD;
    SS15[27][24] = 4'hC;
    SS15[28][24] = 4'hC;
    SS15[29][24] = 4'hC;
    SS15[30][24] = 4'hD;
    SS15[31][24] = 4'hD;
    SS15[32][24] = 4'hD;
    SS15[33][24] = 4'h3;
    SS15[34][24] = 4'h3;
    SS15[35][24] = 4'h3;
    SS15[36][24] = 4'h3;
    SS15[37][24] = 4'h0;
    SS15[38][24] = 4'h0;
    SS15[39][24] = 4'h0;
    SS15[40][24] = 4'h0;
    SS15[41][24] = 4'h0;
    SS15[42][24] = 4'h0;
    SS15[43][24] = 4'h0;
    SS15[44][24] = 4'h0;
    SS15[45][24] = 4'h0;
    SS15[46][24] = 4'h0;
    SS15[47][24] = 4'h0;
    SS15[0][25] = 4'h0;
    SS15[1][25] = 4'h0;
    SS15[2][25] = 4'h0;
    SS15[3][25] = 4'h0;
    SS15[4][25] = 4'hE;
    SS15[5][25] = 4'hE;
    SS15[6][25] = 4'hE;
    SS15[7][25] = 4'hE;
    SS15[8][25] = 4'hE;
    SS15[9][25] = 4'hE;
    SS15[10][25] = 4'hE;
    SS15[11][25] = 4'hC;
    SS15[12][25] = 4'hE;
    SS15[13][25] = 4'hE;
    SS15[14][25] = 4'hC;
    SS15[15][25] = 4'hC;
    SS15[16][25] = 4'hC;
    SS15[17][25] = 4'hC;
    SS15[18][25] = 4'hC;
    SS15[19][25] = 4'hC;
    SS15[20][25] = 4'hC;
    SS15[21][25] = 4'hC;
    SS15[22][25] = 4'hC;
    SS15[23][25] = 4'hC;
    SS15[24][25] = 4'hC;
    SS15[25][25] = 4'hC;
    SS15[26][25] = 4'hC;
    SS15[27][25] = 4'hC;
    SS15[28][25] = 4'hC;
    SS15[29][25] = 4'hC;
    SS15[30][25] = 4'hD;
    SS15[31][25] = 4'hD;
    SS15[32][25] = 4'hD;
    SS15[33][25] = 4'hD;
    SS15[34][25] = 4'hD;
    SS15[35][25] = 4'h3;
    SS15[36][25] = 4'h0;
    SS15[37][25] = 4'h0;
    SS15[38][25] = 4'h0;
    SS15[39][25] = 4'h0;
    SS15[40][25] = 4'h0;
    SS15[41][25] = 4'h0;
    SS15[42][25] = 4'h0;
    SS15[43][25] = 4'h0;
    SS15[44][25] = 4'h0;
    SS15[45][25] = 4'h0;
    SS15[46][25] = 4'h0;
    SS15[47][25] = 4'h0;
    SS15[0][26] = 4'h0;
    SS15[1][26] = 4'h0;
    SS15[2][26] = 4'h0;
    SS15[3][26] = 4'h0;
    SS15[4][26] = 4'h0;
    SS15[5][26] = 4'h0;
    SS15[6][26] = 4'h0;
    SS15[7][26] = 4'hE;
    SS15[8][26] = 4'hE;
    SS15[9][26] = 4'hE;
    SS15[10][26] = 4'hC;
    SS15[11][26] = 4'hC;
    SS15[12][26] = 4'hC;
    SS15[13][26] = 4'hC;
    SS15[14][26] = 4'hC;
    SS15[15][26] = 4'hC;
    SS15[16][26] = 4'hC;
    SS15[17][26] = 4'hC;
    SS15[18][26] = 4'hC;
    SS15[19][26] = 4'hC;
    SS15[20][26] = 4'hD;
    SS15[21][26] = 4'hD;
    SS15[22][26] = 4'hC;
    SS15[23][26] = 4'hC;
    SS15[24][26] = 4'hC;
    SS15[25][26] = 4'hC;
    SS15[26][26] = 4'hC;
    SS15[27][26] = 4'hC;
    SS15[28][26] = 4'hC;
    SS15[29][26] = 4'hE;
    SS15[30][26] = 4'hD;
    SS15[31][26] = 4'hD;
    SS15[32][26] = 4'hD;
    SS15[33][26] = 4'hD;
    SS15[34][26] = 4'hD;
    SS15[35][26] = 4'hD;
    SS15[36][26] = 4'h0;
    SS15[37][26] = 4'h0;
    SS15[38][26] = 4'h0;
    SS15[39][26] = 4'h0;
    SS15[40][26] = 4'h0;
    SS15[41][26] = 4'h0;
    SS15[42][26] = 4'h0;
    SS15[43][26] = 4'h0;
    SS15[44][26] = 4'h0;
    SS15[45][26] = 4'h0;
    SS15[46][26] = 4'h0;
    SS15[47][26] = 4'h0;
    SS15[0][27] = 4'h0;
    SS15[1][27] = 4'h0;
    SS15[2][27] = 4'h0;
    SS15[3][27] = 4'h0;
    SS15[4][27] = 4'h0;
    SS15[5][27] = 4'h0;
    SS15[6][27] = 4'h0;
    SS15[7][27] = 4'h0;
    SS15[8][27] = 4'h0;
    SS15[9][27] = 4'hE;
    SS15[10][27] = 4'hC;
    SS15[11][27] = 4'hC;
    SS15[12][27] = 4'hC;
    SS15[13][27] = 4'hC;
    SS15[14][27] = 4'hC;
    SS15[15][27] = 4'hC;
    SS15[16][27] = 4'hC;
    SS15[17][27] = 4'hC;
    SS15[18][27] = 4'hC;
    SS15[19][27] = 4'hD;
    SS15[20][27] = 4'hD;
    SS15[21][27] = 4'hD;
    SS15[22][27] = 4'hD;
    SS15[23][27] = 4'hD;
    SS15[24][27] = 4'hD;
    SS15[25][27] = 4'hC;
    SS15[26][27] = 4'hC;
    SS15[27][27] = 4'hC;
    SS15[28][27] = 4'hC;
    SS15[29][27] = 4'hE;
    SS15[30][27] = 4'hE;
    SS15[31][27] = 4'hE;
    SS15[32][27] = 4'hD;
    SS15[33][27] = 4'hD;
    SS15[34][27] = 4'hD;
    SS15[35][27] = 4'h0;
    SS15[36][27] = 4'h0;
    SS15[37][27] = 4'h0;
    SS15[38][27] = 4'h0;
    SS15[39][27] = 4'h0;
    SS15[40][27] = 4'h0;
    SS15[41][27] = 4'h0;
    SS15[42][27] = 4'h0;
    SS15[43][27] = 4'h0;
    SS15[44][27] = 4'h0;
    SS15[45][27] = 4'h0;
    SS15[46][27] = 4'h0;
    SS15[47][27] = 4'h0;
    SS15[0][28] = 4'h0;
    SS15[1][28] = 4'h0;
    SS15[2][28] = 4'h0;
    SS15[3][28] = 4'h0;
    SS15[4][28] = 4'h0;
    SS15[5][28] = 4'h0;
    SS15[6][28] = 4'h0;
    SS15[7][28] = 4'h0;
    SS15[8][28] = 4'h0;
    SS15[9][28] = 4'hC;
    SS15[10][28] = 4'hC;
    SS15[11][28] = 4'hC;
    SS15[12][28] = 4'hC;
    SS15[13][28] = 4'hC;
    SS15[14][28] = 4'hC;
    SS15[15][28] = 4'hC;
    SS15[16][28] = 4'hC;
    SS15[17][28] = 4'hC;
    SS15[18][28] = 4'hC;
    SS15[19][28] = 4'hD;
    SS15[20][28] = 4'hD;
    SS15[21][28] = 4'hD;
    SS15[22][28] = 4'hD;
    SS15[23][28] = 4'hD;
    SS15[24][28] = 4'hD;
    SS15[25][28] = 4'hC;
    SS15[26][28] = 4'hC;
    SS15[27][28] = 4'hC;
    SS15[28][28] = 4'hC;
    SS15[29][28] = 4'hE;
    SS15[30][28] = 4'hE;
    SS15[31][28] = 4'hE;
    SS15[32][28] = 4'hD;
    SS15[33][28] = 4'hD;
    SS15[34][28] = 4'hD;
    SS15[35][28] = 4'h0;
    SS15[36][28] = 4'h0;
    SS15[37][28] = 4'h0;
    SS15[38][28] = 4'h0;
    SS15[39][28] = 4'h0;
    SS15[40][28] = 4'h0;
    SS15[41][28] = 4'h0;
    SS15[42][28] = 4'h0;
    SS15[43][28] = 4'h0;
    SS15[44][28] = 4'h0;
    SS15[45][28] = 4'h0;
    SS15[46][28] = 4'h0;
    SS15[47][28] = 4'h0;
    SS15[0][29] = 4'h0;
    SS15[1][29] = 4'h0;
    SS15[2][29] = 4'h0;
    SS15[3][29] = 4'h0;
    SS15[4][29] = 4'h0;
    SS15[5][29] = 4'h0;
    SS15[6][29] = 4'h0;
    SS15[7][29] = 4'h0;
    SS15[8][29] = 4'h0;
    SS15[9][29] = 4'hC;
    SS15[10][29] = 4'hC;
    SS15[11][29] = 4'hC;
    SS15[12][29] = 4'hC;
    SS15[13][29] = 4'hC;
    SS15[14][29] = 4'hC;
    SS15[15][29] = 4'hC;
    SS15[16][29] = 4'hC;
    SS15[17][29] = 4'hC;
    SS15[18][29] = 4'hC;
    SS15[19][29] = 4'hE;
    SS15[20][29] = 4'hE;
    SS15[21][29] = 4'hE;
    SS15[22][29] = 4'hD;
    SS15[23][29] = 4'hD;
    SS15[24][29] = 4'hD;
    SS15[25][29] = 4'hC;
    SS15[26][29] = 4'hC;
    SS15[27][29] = 4'hC;
    SS15[28][29] = 4'hC;
    SS15[29][29] = 4'hC;
    SS15[30][29] = 4'hE;
    SS15[31][29] = 4'hD;
    SS15[32][29] = 4'hD;
    SS15[33][29] = 4'hD;
    SS15[34][29] = 4'hD;
    SS15[35][29] = 4'hD;
    SS15[36][29] = 4'hD;
    SS15[37][29] = 4'h0;
    SS15[38][29] = 4'h0;
    SS15[39][29] = 4'h0;
    SS15[40][29] = 4'h0;
    SS15[41][29] = 4'h0;
    SS15[42][29] = 4'h0;
    SS15[43][29] = 4'h0;
    SS15[44][29] = 4'h0;
    SS15[45][29] = 4'h0;
    SS15[46][29] = 4'h0;
    SS15[47][29] = 4'h0;
    SS15[0][30] = 4'h0;
    SS15[1][30] = 4'h0;
    SS15[2][30] = 4'h0;
    SS15[3][30] = 4'h0;
    SS15[4][30] = 4'h0;
    SS15[5][30] = 4'h0;
    SS15[6][30] = 4'h0;
    SS15[7][30] = 4'h0;
    SS15[8][30] = 4'hC;
    SS15[9][30] = 4'hC;
    SS15[10][30] = 4'hC;
    SS15[11][30] = 4'hC;
    SS15[12][30] = 4'hC;
    SS15[13][30] = 4'hC;
    SS15[14][30] = 4'hC;
    SS15[15][30] = 4'hD;
    SS15[16][30] = 4'hC;
    SS15[17][30] = 4'hC;
    SS15[18][30] = 4'hE;
    SS15[19][30] = 4'hE;
    SS15[20][30] = 4'hE;
    SS15[21][30] = 4'hE;
    SS15[22][30] = 4'hE;
    SS15[23][30] = 4'hE;
    SS15[24][30] = 4'hD;
    SS15[25][30] = 4'hC;
    SS15[26][30] = 4'hC;
    SS15[27][30] = 4'hC;
    SS15[28][30] = 4'hC;
    SS15[29][30] = 4'hC;
    SS15[30][30] = 4'hC;
    SS15[31][30] = 4'hE;
    SS15[32][30] = 4'hD;
    SS15[33][30] = 4'hD;
    SS15[34][30] = 4'hD;
    SS15[35][30] = 4'hD;
    SS15[36][30] = 4'hD;
    SS15[37][30] = 4'h3;
    SS15[38][30] = 4'h3;
    SS15[39][30] = 4'h3;
    SS15[40][30] = 4'h0;
    SS15[41][30] = 4'h0;
    SS15[42][30] = 4'h0;
    SS15[43][30] = 4'h0;
    SS15[44][30] = 4'h0;
    SS15[45][30] = 4'h0;
    SS15[46][30] = 4'h0;
    SS15[47][30] = 4'h0;
    SS15[0][31] = 4'h0;
    SS15[1][31] = 4'h0;
    SS15[2][31] = 4'h0;
    SS15[3][31] = 4'h0;
    SS15[4][31] = 4'h0;
    SS15[5][31] = 4'h0;
    SS15[6][31] = 4'h0;
    SS15[7][31] = 4'h0;
    SS15[8][31] = 4'hC;
    SS15[9][31] = 4'hC;
    SS15[10][31] = 4'hC;
    SS15[11][31] = 4'hC;
    SS15[12][31] = 4'hC;
    SS15[13][31] = 4'hC;
    SS15[14][31] = 4'hD;
    SS15[15][31] = 4'hD;
    SS15[16][31] = 4'hD;
    SS15[17][31] = 4'hD;
    SS15[18][31] = 4'hE;
    SS15[19][31] = 4'hE;
    SS15[20][31] = 4'hE;
    SS15[21][31] = 4'hE;
    SS15[22][31] = 4'hE;
    SS15[23][31] = 4'hE;
    SS15[24][31] = 4'hC;
    SS15[25][31] = 4'hC;
    SS15[26][31] = 4'hC;
    SS15[27][31] = 4'hC;
    SS15[28][31] = 4'hC;
    SS15[29][31] = 4'hC;
    SS15[30][31] = 4'hC;
    SS15[31][31] = 4'hE;
    SS15[32][31] = 4'hE;
    SS15[33][31] = 4'hE;
    SS15[34][31] = 4'hD;
    SS15[35][31] = 4'hD;
    SS15[36][31] = 4'hD;
    SS15[37][31] = 4'h3;
    SS15[38][31] = 4'h3;
    SS15[39][31] = 4'h3;
    SS15[40][31] = 4'h0;
    SS15[41][31] = 4'h0;
    SS15[42][31] = 4'h0;
    SS15[43][31] = 4'h0;
    SS15[44][31] = 4'h0;
    SS15[45][31] = 4'h0;
    SS15[46][31] = 4'h0;
    SS15[47][31] = 4'h0;
    SS15[0][32] = 4'h0;
    SS15[1][32] = 4'h0;
    SS15[2][32] = 4'h0;
    SS15[3][32] = 4'h0;
    SS15[4][32] = 4'hC;
    SS15[5][32] = 4'hC;
    SS15[6][32] = 4'h0;
    SS15[7][32] = 4'h0;
    SS15[8][32] = 4'hC;
    SS15[9][32] = 4'hC;
    SS15[10][32] = 4'hC;
    SS15[11][32] = 4'hD;
    SS15[12][32] = 4'hD;
    SS15[13][32] = 4'hD;
    SS15[14][32] = 4'hD;
    SS15[15][32] = 4'hD;
    SS15[16][32] = 4'hD;
    SS15[17][32] = 4'hE;
    SS15[18][32] = 4'hE;
    SS15[19][32] = 4'hE;
    SS15[20][32] = 4'hE;
    SS15[21][32] = 4'hE;
    SS15[22][32] = 4'hE;
    SS15[23][32] = 4'hE;
    SS15[24][32] = 4'hC;
    SS15[25][32] = 4'hC;
    SS15[26][32] = 4'hC;
    SS15[27][32] = 4'hC;
    SS15[28][32] = 4'hC;
    SS15[29][32] = 4'hC;
    SS15[30][32] = 4'hE;
    SS15[31][32] = 4'hE;
    SS15[32][32] = 4'hE;
    SS15[33][32] = 4'hE;
    SS15[34][32] = 4'hE;
    SS15[35][32] = 4'hE;
    SS15[36][32] = 4'hE;
    SS15[37][32] = 4'h3;
    SS15[38][32] = 4'h3;
    SS15[39][32] = 4'h3;
    SS15[40][32] = 4'h0;
    SS15[41][32] = 4'h0;
    SS15[42][32] = 4'h0;
    SS15[43][32] = 4'h0;
    SS15[44][32] = 4'h0;
    SS15[45][32] = 4'h0;
    SS15[46][32] = 4'h0;
    SS15[47][32] = 4'h0;
    SS15[0][33] = 4'h0;
    SS15[1][33] = 4'h0;
    SS15[2][33] = 4'h0;
    SS15[3][33] = 4'h0;
    SS15[4][33] = 4'hC;
    SS15[5][33] = 4'hC;
    SS15[6][33] = 4'hC;
    SS15[7][33] = 4'hC;
    SS15[8][33] = 4'hC;
    SS15[9][33] = 4'hC;
    SS15[10][33] = 4'hD;
    SS15[11][33] = 4'hD;
    SS15[12][33] = 4'hD;
    SS15[13][33] = 4'hD;
    SS15[14][33] = 4'hE;
    SS15[15][33] = 4'hE;
    SS15[16][33] = 4'hD;
    SS15[17][33] = 4'hE;
    SS15[18][33] = 4'hE;
    SS15[19][33] = 4'hE;
    SS15[20][33] = 4'hE;
    SS15[21][33] = 4'hE;
    SS15[22][33] = 4'hE;
    SS15[23][33] = 4'hD;
    SS15[24][33] = 4'hC;
    SS15[25][33] = 4'hC;
    SS15[26][33] = 4'hC;
    SS15[27][33] = 4'hC;
    SS15[28][33] = 4'hC;
    SS15[29][33] = 4'hC;
    SS15[30][33] = 4'hC;
    SS15[31][33] = 4'hE;
    SS15[32][33] = 4'hE;
    SS15[33][33] = 4'hE;
    SS15[34][33] = 4'hE;
    SS15[35][33] = 4'hE;
    SS15[36][33] = 4'hD;
    SS15[37][33] = 4'hD;
    SS15[38][33] = 4'hD;
    SS15[39][33] = 4'h0;
    SS15[40][33] = 4'h0;
    SS15[41][33] = 4'h0;
    SS15[42][33] = 4'h0;
    SS15[43][33] = 4'h0;
    SS15[44][33] = 4'h0;
    SS15[45][33] = 4'h0;
    SS15[46][33] = 4'h0;
    SS15[47][33] = 4'h0;
    SS15[0][34] = 4'h0;
    SS15[1][34] = 4'h0;
    SS15[2][34] = 4'h0;
    SS15[3][34] = 4'h0;
    SS15[4][34] = 4'hC;
    SS15[5][34] = 4'hC;
    SS15[6][34] = 4'hC;
    SS15[7][34] = 4'hC;
    SS15[8][34] = 4'hC;
    SS15[9][34] = 4'hC;
    SS15[10][34] = 4'hE;
    SS15[11][34] = 4'hD;
    SS15[12][34] = 4'hD;
    SS15[13][34] = 4'hE;
    SS15[14][34] = 4'hE;
    SS15[15][34] = 4'hE;
    SS15[16][34] = 4'h0;
    SS15[17][34] = 4'h0;
    SS15[18][34] = 4'hE;
    SS15[19][34] = 4'hE;
    SS15[20][34] = 4'hE;
    SS15[21][34] = 4'hE;
    SS15[22][34] = 4'hE;
    SS15[23][34] = 4'hD;
    SS15[24][34] = 4'hD;
    SS15[25][34] = 4'hD;
    SS15[26][34] = 4'hC;
    SS15[27][34] = 4'hC;
    SS15[28][34] = 4'hC;
    SS15[29][34] = 4'hC;
    SS15[30][34] = 4'hC;
    SS15[31][34] = 4'hC;
    SS15[32][34] = 4'hE;
    SS15[33][34] = 4'hE;
    SS15[34][34] = 4'hE;
    SS15[35][34] = 4'hE;
    SS15[36][34] = 4'hD;
    SS15[37][34] = 4'hD;
    SS15[38][34] = 4'hD;
    SS15[39][34] = 4'hD;
    SS15[40][34] = 4'hD;
    SS15[41][34] = 4'hD;
    SS15[42][34] = 4'h0;
    SS15[43][34] = 4'h0;
    SS15[44][34] = 4'h0;
    SS15[45][34] = 4'h0;
    SS15[46][34] = 4'h0;
    SS15[47][34] = 4'h0;
    SS15[0][35] = 4'h0;
    SS15[1][35] = 4'h0;
    SS15[2][35] = 4'h0;
    SS15[3][35] = 4'hC;
    SS15[4][35] = 4'hC;
    SS15[5][35] = 4'hC;
    SS15[6][35] = 4'hC;
    SS15[7][35] = 4'hC;
    SS15[8][35] = 4'hC;
    SS15[9][35] = 4'hC;
    SS15[10][35] = 4'hE;
    SS15[11][35] = 4'hE;
    SS15[12][35] = 4'hE;
    SS15[13][35] = 4'hE;
    SS15[14][35] = 4'hE;
    SS15[15][35] = 4'hE;
    SS15[16][35] = 4'h0;
    SS15[17][35] = 4'h0;
    SS15[18][35] = 4'h0;
    SS15[19][35] = 4'h0;
    SS15[20][35] = 4'h0;
    SS15[21][35] = 4'hE;
    SS15[22][35] = 4'hD;
    SS15[23][35] = 4'hD;
    SS15[24][35] = 4'hD;
    SS15[25][35] = 4'hD;
    SS15[26][35] = 4'hC;
    SS15[27][35] = 4'hC;
    SS15[28][35] = 4'hC;
    SS15[29][35] = 4'hC;
    SS15[30][35] = 4'hC;
    SS15[31][35] = 4'hC;
    SS15[32][35] = 4'hE;
    SS15[33][35] = 4'hE;
    SS15[34][35] = 4'hE;
    SS15[35][35] = 4'hE;
    SS15[36][35] = 4'hD;
    SS15[37][35] = 4'hD;
    SS15[38][35] = 4'hD;
    SS15[39][35] = 4'hD;
    SS15[40][35] = 4'hD;
    SS15[41][35] = 4'hD;
    SS15[42][35] = 4'h0;
    SS15[43][35] = 4'h0;
    SS15[44][35] = 4'h0;
    SS15[45][35] = 4'h0;
    SS15[46][35] = 4'h0;
    SS15[47][35] = 4'h0;
    SS15[0][36] = 4'h0;
    SS15[1][36] = 4'h0;
    SS15[2][36] = 4'h0;
    SS15[3][36] = 4'hC;
    SS15[4][36] = 4'hC;
    SS15[5][36] = 4'hC;
    SS15[6][36] = 4'hD;
    SS15[7][36] = 4'hD;
    SS15[8][36] = 4'hC;
    SS15[9][36] = 4'hE;
    SS15[10][36] = 4'hE;
    SS15[11][36] = 4'hE;
    SS15[12][36] = 4'h0;
    SS15[13][36] = 4'h0;
    SS15[14][36] = 4'h0;
    SS15[15][36] = 4'hE;
    SS15[16][36] = 4'h0;
    SS15[17][36] = 4'h0;
    SS15[18][36] = 4'h0;
    SS15[19][36] = 4'h0;
    SS15[20][36] = 4'h0;
    SS15[21][36] = 4'h0;
    SS15[22][36] = 4'hE;
    SS15[23][36] = 4'hD;
    SS15[24][36] = 4'hD;
    SS15[25][36] = 4'hC;
    SS15[26][36] = 4'hC;
    SS15[27][36] = 4'hC;
    SS15[28][36] = 4'hC;
    SS15[29][36] = 4'hC;
    SS15[30][36] = 4'hC;
    SS15[31][36] = 4'hC;
    SS15[32][36] = 4'hE;
    SS15[33][36] = 4'hE;
    SS15[34][36] = 4'hE;
    SS15[35][36] = 4'hE;
    SS15[36][36] = 4'hE;
    SS15[37][36] = 4'hE;
    SS15[38][36] = 4'hD;
    SS15[39][36] = 4'hD;
    SS15[40][36] = 4'hD;
    SS15[41][36] = 4'h0;
    SS15[42][36] = 4'h0;
    SS15[43][36] = 4'h0;
    SS15[44][36] = 4'h0;
    SS15[45][36] = 4'h0;
    SS15[46][36] = 4'h0;
    SS15[47][36] = 4'h0;
    SS15[0][37] = 4'h0;
    SS15[1][37] = 4'h0;
    SS15[2][37] = 4'hC;
    SS15[3][37] = 4'hC;
    SS15[4][37] = 4'hC;
    SS15[5][37] = 4'hC;
    SS15[6][37] = 4'hD;
    SS15[7][37] = 4'hD;
    SS15[8][37] = 4'hD;
    SS15[9][37] = 4'h0;
    SS15[10][37] = 4'hE;
    SS15[11][37] = 4'hE;
    SS15[12][37] = 4'h0;
    SS15[13][37] = 4'h0;
    SS15[14][37] = 4'h0;
    SS15[15][37] = 4'h0;
    SS15[16][37] = 4'h0;
    SS15[17][37] = 4'h0;
    SS15[18][37] = 4'h0;
    SS15[19][37] = 4'h0;
    SS15[20][37] = 4'h0;
    SS15[21][37] = 4'h0;
    SS15[22][37] = 4'hE;
    SS15[23][37] = 4'hE;
    SS15[24][37] = 4'hE;
    SS15[25][37] = 4'hD;
    SS15[26][37] = 4'hC;
    SS15[27][37] = 4'hC;
    SS15[28][37] = 4'hC;
    SS15[29][37] = 4'hC;
    SS15[30][37] = 4'hC;
    SS15[31][37] = 4'h0;
    SS15[32][37] = 4'h0;
    SS15[33][37] = 4'hE;
    SS15[34][37] = 4'hE;
    SS15[35][37] = 4'hE;
    SS15[36][37] = 4'hE;
    SS15[37][37] = 4'hE;
    SS15[38][37] = 4'hD;
    SS15[39][37] = 4'hD;
    SS15[40][37] = 4'hD;
    SS15[41][37] = 4'h0;
    SS15[42][37] = 4'h0;
    SS15[43][37] = 4'h0;
    SS15[44][37] = 4'h0;
    SS15[45][37] = 4'h0;
    SS15[46][37] = 4'h0;
    SS15[47][37] = 4'h0;
    SS15[0][38] = 4'h0;
    SS15[1][38] = 4'h0;
    SS15[2][38] = 4'hD;
    SS15[3][38] = 4'hD;
    SS15[4][38] = 4'hD;
    SS15[5][38] = 4'hD;
    SS15[6][38] = 4'hD;
    SS15[7][38] = 4'hD;
    SS15[8][38] = 4'h0;
    SS15[9][38] = 4'h0;
    SS15[10][38] = 4'h0;
    SS15[11][38] = 4'h0;
    SS15[12][38] = 4'h0;
    SS15[13][38] = 4'h0;
    SS15[14][38] = 4'h0;
    SS15[15][38] = 4'h0;
    SS15[16][38] = 4'h0;
    SS15[17][38] = 4'h0;
    SS15[18][38] = 4'h0;
    SS15[19][38] = 4'h0;
    SS15[20][38] = 4'h0;
    SS15[21][38] = 4'hE;
    SS15[22][38] = 4'hE;
    SS15[23][38] = 4'hE;
    SS15[24][38] = 4'hD;
    SS15[25][38] = 4'hD;
    SS15[26][38] = 4'hD;
    SS15[27][38] = 4'hD;
    SS15[28][38] = 4'hC;
    SS15[29][38] = 4'hC;
    SS15[30][38] = 4'hC;
    SS15[31][38] = 4'h0;
    SS15[32][38] = 4'h0;
    SS15[33][38] = 4'h0;
    SS15[34][38] = 4'h0;
    SS15[35][38] = 4'h0;
    SS15[36][38] = 4'hE;
    SS15[37][38] = 4'hD;
    SS15[38][38] = 4'hD;
    SS15[39][38] = 4'hD;
    SS15[40][38] = 4'hD;
    SS15[41][38] = 4'hD;
    SS15[42][38] = 4'hD;
    SS15[43][38] = 4'hD;
    SS15[44][38] = 4'h0;
    SS15[45][38] = 4'h0;
    SS15[46][38] = 4'h0;
    SS15[47][38] = 4'h0;
    SS15[0][39] = 4'h0;
    SS15[1][39] = 4'h0;
    SS15[2][39] = 4'hD;
    SS15[3][39] = 4'hD;
    SS15[4][39] = 4'hD;
    SS15[5][39] = 4'h0;
    SS15[6][39] = 4'h0;
    SS15[7][39] = 4'hD;
    SS15[8][39] = 4'h0;
    SS15[9][39] = 4'h0;
    SS15[10][39] = 4'h0;
    SS15[11][39] = 4'h0;
    SS15[12][39] = 4'h0;
    SS15[13][39] = 4'h0;
    SS15[14][39] = 4'h0;
    SS15[15][39] = 4'h0;
    SS15[16][39] = 4'h0;
    SS15[17][39] = 4'h0;
    SS15[18][39] = 4'h0;
    SS15[19][39] = 4'h0;
    SS15[20][39] = 4'h0;
    SS15[21][39] = 4'h0;
    SS15[22][39] = 4'h0;
    SS15[23][39] = 4'hE;
    SS15[24][39] = 4'hD;
    SS15[25][39] = 4'hD;
    SS15[26][39] = 4'hD;
    SS15[27][39] = 4'hC;
    SS15[28][39] = 4'hC;
    SS15[29][39] = 4'hC;
    SS15[30][39] = 4'h0;
    SS15[31][39] = 4'h0;
    SS15[32][39] = 4'h0;
    SS15[33][39] = 4'h0;
    SS15[34][39] = 4'h0;
    SS15[35][39] = 4'h0;
    SS15[36][39] = 4'h0;
    SS15[37][39] = 4'h0;
    SS15[38][39] = 4'hD;
    SS15[39][39] = 4'hD;
    SS15[40][39] = 4'hD;
    SS15[41][39] = 4'hD;
    SS15[42][39] = 4'hD;
    SS15[43][39] = 4'h0;
    SS15[44][39] = 4'h0;
    SS15[45][39] = 4'h0;
    SS15[46][39] = 4'h0;
    SS15[47][39] = 4'h0;
    SS15[0][40] = 4'h0;
    SS15[1][40] = 4'h0;
    SS15[2][40] = 4'hD;
    SS15[3][40] = 4'hD;
    SS15[4][40] = 4'h0;
    SS15[5][40] = 4'h0;
    SS15[6][40] = 4'h0;
    SS15[7][40] = 4'h0;
    SS15[8][40] = 4'h0;
    SS15[9][40] = 4'h0;
    SS15[10][40] = 4'h0;
    SS15[11][40] = 4'h0;
    SS15[12][40] = 4'h0;
    SS15[13][40] = 4'h0;
    SS15[14][40] = 4'h0;
    SS15[15][40] = 4'h0;
    SS15[16][40] = 4'h0;
    SS15[17][40] = 4'h0;
    SS15[18][40] = 4'h0;
    SS15[19][40] = 4'h0;
    SS15[20][40] = 4'h0;
    SS15[21][40] = 4'h0;
    SS15[22][40] = 4'h0;
    SS15[23][40] = 4'h0;
    SS15[24][40] = 4'hE;
    SS15[25][40] = 4'hD;
    SS15[26][40] = 4'hD;
    SS15[27][40] = 4'hC;
    SS15[28][40] = 4'hC;
    SS15[29][40] = 4'hC;
    SS15[30][40] = 4'h0;
    SS15[31][40] = 4'h0;
    SS15[32][40] = 4'h0;
    SS15[33][40] = 4'h0;
    SS15[34][40] = 4'h0;
    SS15[35][40] = 4'h0;
    SS15[36][40] = 4'h0;
    SS15[37][40] = 4'h0;
    SS15[38][40] = 4'h0;
    SS15[39][40] = 4'h0;
    SS15[40][40] = 4'h0;
    SS15[41][40] = 4'hD;
    SS15[42][40] = 4'hD;
    SS15[43][40] = 4'h0;
    SS15[44][40] = 4'h0;
    SS15[45][40] = 4'h0;
    SS15[46][40] = 4'h0;
    SS15[47][40] = 4'h0;
    SS15[0][41] = 4'h0;
    SS15[1][41] = 4'h0;
    SS15[2][41] = 4'h0;
    SS15[3][41] = 4'h0;
    SS15[4][41] = 4'h0;
    SS15[5][41] = 4'h0;
    SS15[6][41] = 4'h0;
    SS15[7][41] = 4'h0;
    SS15[8][41] = 4'h0;
    SS15[9][41] = 4'h0;
    SS15[10][41] = 4'h0;
    SS15[11][41] = 4'h0;
    SS15[12][41] = 4'h0;
    SS15[13][41] = 4'h0;
    SS15[14][41] = 4'h0;
    SS15[15][41] = 4'h0;
    SS15[16][41] = 4'h0;
    SS15[17][41] = 4'h0;
    SS15[18][41] = 4'h0;
    SS15[19][41] = 4'h0;
    SS15[20][41] = 4'h0;
    SS15[21][41] = 4'h0;
    SS15[22][41] = 4'h0;
    SS15[23][41] = 4'hE;
    SS15[24][41] = 4'hE;
    SS15[25][41] = 4'hE;
    SS15[26][41] = 4'hC;
    SS15[27][41] = 4'hC;
    SS15[28][41] = 4'hC;
    SS15[29][41] = 4'hC;
    SS15[30][41] = 4'h0;
    SS15[31][41] = 4'h0;
    SS15[32][41] = 4'h0;
    SS15[33][41] = 4'h0;
    SS15[34][41] = 4'h0;
    SS15[35][41] = 4'h0;
    SS15[36][41] = 4'h0;
    SS15[37][41] = 4'h0;
    SS15[38][41] = 4'h0;
    SS15[39][41] = 4'h0;
    SS15[40][41] = 4'h0;
    SS15[41][41] = 4'h0;
    SS15[42][41] = 4'h0;
    SS15[43][41] = 4'h0;
    SS15[44][41] = 4'h0;
    SS15[45][41] = 4'h0;
    SS15[46][41] = 4'h0;
    SS15[47][41] = 4'h0;
    SS15[0][42] = 4'h0;
    SS15[1][42] = 4'h0;
    SS15[2][42] = 4'h0;
    SS15[3][42] = 4'h0;
    SS15[4][42] = 4'h0;
    SS15[5][42] = 4'h0;
    SS15[6][42] = 4'h0;
    SS15[7][42] = 4'h0;
    SS15[8][42] = 4'h0;
    SS15[9][42] = 4'h0;
    SS15[10][42] = 4'h0;
    SS15[11][42] = 4'h0;
    SS15[12][42] = 4'h0;
    SS15[13][42] = 4'h0;
    SS15[14][42] = 4'h0;
    SS15[15][42] = 4'h0;
    SS15[16][42] = 4'h0;
    SS15[17][42] = 4'h0;
    SS15[18][42] = 4'h0;
    SS15[19][42] = 4'h0;
    SS15[20][42] = 4'h0;
    SS15[21][42] = 4'h0;
    SS15[22][42] = 4'h0;
    SS15[23][42] = 4'hE;
    SS15[24][42] = 4'hE;
    SS15[25][42] = 4'hE;
    SS15[26][42] = 4'hC;
    SS15[27][42] = 4'hC;
    SS15[28][42] = 4'hC;
    SS15[29][42] = 4'hC;
    SS15[30][42] = 4'h0;
    SS15[31][42] = 4'h0;
    SS15[32][42] = 4'h0;
    SS15[33][42] = 4'h0;
    SS15[34][42] = 4'h0;
    SS15[35][42] = 4'h0;
    SS15[36][42] = 4'h0;
    SS15[37][42] = 4'h0;
    SS15[38][42] = 4'h0;
    SS15[39][42] = 4'h0;
    SS15[40][42] = 4'h0;
    SS15[41][42] = 4'h0;
    SS15[42][42] = 4'h0;
    SS15[43][42] = 4'h0;
    SS15[44][42] = 4'h0;
    SS15[45][42] = 4'h0;
    SS15[46][42] = 4'h0;
    SS15[47][42] = 4'h0;
    SS15[0][43] = 4'h0;
    SS15[1][43] = 4'h0;
    SS15[2][43] = 4'h0;
    SS15[3][43] = 4'h0;
    SS15[4][43] = 4'h0;
    SS15[5][43] = 4'h0;
    SS15[6][43] = 4'h0;
    SS15[7][43] = 4'h0;
    SS15[8][43] = 4'h0;
    SS15[9][43] = 4'h0;
    SS15[10][43] = 4'h0;
    SS15[11][43] = 4'h0;
    SS15[12][43] = 4'h0;
    SS15[13][43] = 4'h0;
    SS15[14][43] = 4'h0;
    SS15[15][43] = 4'h0;
    SS15[16][43] = 4'h0;
    SS15[17][43] = 4'h0;
    SS15[18][43] = 4'h0;
    SS15[19][43] = 4'h0;
    SS15[20][43] = 4'h0;
    SS15[21][43] = 4'h0;
    SS15[22][43] = 4'h0;
    SS15[23][43] = 4'h0;
    SS15[24][43] = 4'h0;
    SS15[25][43] = 4'hE;
    SS15[26][43] = 4'hC;
    SS15[27][43] = 4'hC;
    SS15[28][43] = 4'hC;
    SS15[29][43] = 4'hC;
    SS15[30][43] = 4'hC;
    SS15[31][43] = 4'hC;
    SS15[32][43] = 4'h0;
    SS15[33][43] = 4'h0;
    SS15[34][43] = 4'h0;
    SS15[35][43] = 4'h0;
    SS15[36][43] = 4'h0;
    SS15[37][43] = 4'h0;
    SS15[38][43] = 4'h0;
    SS15[39][43] = 4'h0;
    SS15[40][43] = 4'h0;
    SS15[41][43] = 4'h0;
    SS15[42][43] = 4'h0;
    SS15[43][43] = 4'h0;
    SS15[44][43] = 4'h0;
    SS15[45][43] = 4'h0;
    SS15[46][43] = 4'h0;
    SS15[47][43] = 4'h0;
    SS15[0][44] = 4'h0;
    SS15[1][44] = 4'h0;
    SS15[2][44] = 4'h0;
    SS15[3][44] = 4'h0;
    SS15[4][44] = 4'h0;
    SS15[5][44] = 4'h0;
    SS15[6][44] = 4'h0;
    SS15[7][44] = 4'h0;
    SS15[8][44] = 4'h0;
    SS15[9][44] = 4'h0;
    SS15[10][44] = 4'h0;
    SS15[11][44] = 4'h0;
    SS15[12][44] = 4'h0;
    SS15[13][44] = 4'h0;
    SS15[14][44] = 4'h0;
    SS15[15][44] = 4'h0;
    SS15[16][44] = 4'h0;
    SS15[17][44] = 4'h0;
    SS15[18][44] = 4'h0;
    SS15[19][44] = 4'h0;
    SS15[20][44] = 4'h0;
    SS15[21][44] = 4'h0;
    SS15[22][44] = 4'h0;
    SS15[23][44] = 4'h0;
    SS15[24][44] = 4'h0;
    SS15[25][44] = 4'hD;
    SS15[26][44] = 4'hD;
    SS15[27][44] = 4'hC;
    SS15[28][44] = 4'hC;
    SS15[29][44] = 4'hC;
    SS15[30][44] = 4'hC;
    SS15[31][44] = 4'hC;
    SS15[32][44] = 4'h0;
    SS15[33][44] = 4'h0;
    SS15[34][44] = 4'h0;
    SS15[35][44] = 4'h0;
    SS15[36][44] = 4'h0;
    SS15[37][44] = 4'h0;
    SS15[38][44] = 4'h0;
    SS15[39][44] = 4'h0;
    SS15[40][44] = 4'h0;
    SS15[41][44] = 4'h0;
    SS15[42][44] = 4'h0;
    SS15[43][44] = 4'h0;
    SS15[44][44] = 4'h0;
    SS15[45][44] = 4'h0;
    SS15[46][44] = 4'h0;
    SS15[47][44] = 4'h0;
    SS15[0][45] = 4'h0;
    SS15[1][45] = 4'h0;
    SS15[2][45] = 4'h0;
    SS15[3][45] = 4'h0;
    SS15[4][45] = 4'h0;
    SS15[5][45] = 4'h0;
    SS15[6][45] = 4'h0;
    SS15[7][45] = 4'h0;
    SS15[8][45] = 4'h0;
    SS15[9][45] = 4'h0;
    SS15[10][45] = 4'h0;
    SS15[11][45] = 4'h0;
    SS15[12][45] = 4'h0;
    SS15[13][45] = 4'h0;
    SS15[14][45] = 4'h0;
    SS15[15][45] = 4'h0;
    SS15[16][45] = 4'h0;
    SS15[17][45] = 4'h0;
    SS15[18][45] = 4'h0;
    SS15[19][45] = 4'h0;
    SS15[20][45] = 4'h0;
    SS15[21][45] = 4'h0;
    SS15[22][45] = 4'h0;
    SS15[23][45] = 4'h0;
    SS15[24][45] = 4'h0;
    SS15[25][45] = 4'hD;
    SS15[26][45] = 4'hD;
    SS15[27][45] = 4'hD;
    SS15[28][45] = 4'hC;
    SS15[29][45] = 4'hC;
    SS15[30][45] = 4'hC;
    SS15[31][45] = 4'h0;
    SS15[32][45] = 4'h0;
    SS15[33][45] = 4'h0;
    SS15[34][45] = 4'h0;
    SS15[35][45] = 4'h0;
    SS15[36][45] = 4'h0;
    SS15[37][45] = 4'h0;
    SS15[38][45] = 4'h0;
    SS15[39][45] = 4'h0;
    SS15[40][45] = 4'h0;
    SS15[41][45] = 4'h0;
    SS15[42][45] = 4'h0;
    SS15[43][45] = 4'h0;
    SS15[44][45] = 4'h0;
    SS15[45][45] = 4'h0;
    SS15[46][45] = 4'h0;
    SS15[47][45] = 4'h0;
    SS15[0][46] = 4'h0;
    SS15[1][46] = 4'h0;
    SS15[2][46] = 4'h0;
    SS15[3][46] = 4'h0;
    SS15[4][46] = 4'h0;
    SS15[5][46] = 4'h0;
    SS15[6][46] = 4'h0;
    SS15[7][46] = 4'h0;
    SS15[8][46] = 4'h0;
    SS15[9][46] = 4'h0;
    SS15[10][46] = 4'h0;
    SS15[11][46] = 4'h0;
    SS15[12][46] = 4'h0;
    SS15[13][46] = 4'h0;
    SS15[14][46] = 4'h0;
    SS15[15][46] = 4'h0;
    SS15[16][46] = 4'h0;
    SS15[17][46] = 4'h0;
    SS15[18][46] = 4'h0;
    SS15[19][46] = 4'h0;
    SS15[20][46] = 4'h0;
    SS15[21][46] = 4'h0;
    SS15[22][46] = 4'h0;
    SS15[23][46] = 4'h0;
    SS15[24][46] = 4'hD;
    SS15[25][46] = 4'hD;
    SS15[26][46] = 4'hD;
    SS15[27][46] = 4'hD;
    SS15[28][46] = 4'hC;
    SS15[29][46] = 4'hC;
    SS15[30][46] = 4'hC;
    SS15[31][46] = 4'h0;
    SS15[32][46] = 4'h0;
    SS15[33][46] = 4'h0;
    SS15[34][46] = 4'h0;
    SS15[35][46] = 4'h0;
    SS15[36][46] = 4'h0;
    SS15[37][46] = 4'h0;
    SS15[38][46] = 4'h0;
    SS15[39][46] = 4'h0;
    SS15[40][46] = 4'h0;
    SS15[41][46] = 4'h0;
    SS15[42][46] = 4'h0;
    SS15[43][46] = 4'h0;
    SS15[44][46] = 4'h0;
    SS15[45][46] = 4'h0;
    SS15[46][46] = 4'h0;
    SS15[47][46] = 4'h0;
    SS15[0][47] = 4'h0;
    SS15[1][47] = 4'h0;
    SS15[2][47] = 4'h0;
    SS15[3][47] = 4'h0;
    SS15[4][47] = 4'h0;
    SS15[5][47] = 4'h0;
    SS15[6][47] = 4'h0;
    SS15[7][47] = 4'h0;
    SS15[8][47] = 4'h0;
    SS15[9][47] = 4'h0;
    SS15[10][47] = 4'h0;
    SS15[11][47] = 4'h0;
    SS15[12][47] = 4'h0;
    SS15[13][47] = 4'h0;
    SS15[14][47] = 4'h0;
    SS15[15][47] = 4'h0;
    SS15[16][47] = 4'h0;
    SS15[17][47] = 4'h0;
    SS15[18][47] = 4'h0;
    SS15[19][47] = 4'h0;
    SS15[20][47] = 4'h0;
    SS15[21][47] = 4'h0;
    SS15[22][47] = 4'h0;
    SS15[23][47] = 4'h0;
    SS15[24][47] = 4'h0;
    SS15[25][47] = 4'h0;
    SS15[26][47] = 4'h0;
    SS15[27][47] = 4'hC;
    SS15[28][47] = 4'hC;
    SS15[29][47] = 4'hC;
    SS15[30][47] = 4'h0;
    SS15[31][47] = 4'h0;
    SS15[32][47] = 4'h0;
    SS15[33][47] = 4'h0;
    SS15[34][47] = 4'h0;
    SS15[35][47] = 4'h0;
    SS15[36][47] = 4'h0;
    SS15[37][47] = 4'h0;
    SS15[38][47] = 4'h0;
    SS15[39][47] = 4'h0;
    SS15[40][47] = 4'h0;
    SS15[41][47] = 4'h0;
    SS15[42][47] = 4'h0;
    SS15[43][47] = 4'h0;
    SS15[44][47] = 4'h0;
    SS15[45][47] = 4'h0;
    SS15[46][47] = 4'h0;
    SS15[47][47] = 4'h0;
 
end
endmodule